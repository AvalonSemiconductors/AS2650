* NGSPICE file created from sid_top.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_4 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_4 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_4 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VNW VPW VSS
.ends

.subckt sid_top DAC_clk DAC_dat_1 DAC_dat_2 DAC_le addr[0] addr[1] addr[2] addr[3]
+ addr[4] addr[5] bus_cyc bus_in[0] bus_in[1] bus_in[2] bus_in[3] bus_in[4] bus_in[5]
+ bus_in[6] bus_in[7] bus_out[0] bus_out[1] bus_out[2] bus_out[3] bus_out[4] bus_out[5]
+ bus_out[6] bus_out[7] bus_we clk rst vdd vss
XFILLER_0_94_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09671_ channels.atk_dec3\[7\] _01991_ _01992_ channels.freq3\[15\] _02055_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_20_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08622_ channels.lfsr\[3\]\[15\] _01122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_171_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13607__A1 _04377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_179_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08553_ channels.clk_div\[0\] _01069_ _01070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_134_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08484_ filters.res_filt\[6\] _01013_ _01014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12830__A2 _04377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09105_ _01554_ _01556_ _01557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__12464__I _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_96_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09036_ _01138_ _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__14335__A2 _05570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12897__A2 _04163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09938_ channels.freq3\[8\] _02248_ _02243_ _02249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10109__B1 channels.ctrl_reg1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13846__A1 _05846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09869_ _02131_ _02194_ _02200_ _00200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_70_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11900_ _03878_ _03879_ _03983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_29_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12880_ _04883_ _04885_ _04886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_158_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11831_ _03891_ _03892_ _03922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12639__I _04644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_116_Left_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14550_ _06544_ _06545_ _06546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_178_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11762_ _03849_ _03851_ _03852_ _03853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_36_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13501_ _05503_ _05506_ _05507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10713_ _02944_ _02969_ _02970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_14481_ _06350_ _06369_ _06478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14854__I _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11693_ _03756_ _03784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_82_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16220_ _08077_ _08092_ _08093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13432_ _05299_ _05358_ _05438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10644_ _02553_ _02575_ _02902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16151_ _07985_ _08001_ _08027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13363_ _05366_ _05368_ _05369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10575_ _02790_ _02829_ _02834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_36_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14790__S _06073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer7 _07362_ net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_114_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_77_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15102_ _07067_ _07068_ _07069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12314_ _03253_ _04224_ _04320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_16082_ _07780_ _07960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_146_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15523__A1 channels.sample3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13294_ _05207_ _05225_ _05300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12337__A1 _03383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15033_ _06958_ _06975_ _07002_ _07003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_20_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12245_ _04234_ _04239_ _04251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_139_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12176_ _04181_ _04182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10899__A1 channels.sample2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11127_ filters.low\[7\] _03345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16984_ _00063_ clknet_leaf_154_clk channels.accum\[0\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15935_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[2\] _07817_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_11058_ _03264_ _03265_ _03266_ _03280_ _00309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_10009_ _02252_ _02291_ _02297_ _00243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_15866_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[2\] _07746_ _07748_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_8_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17605_ _00675_ clknet_leaf_44_clk net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_14817_ filters.band\[20\] _06785_ _06763_ _06803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13065__A2 _05070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15797_ _07693_ _07696_ _00632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17536_ _00606_ clknet_leaf_215_clk channels.exp_periods\[3\]\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14748_ filters.band\[15\] _06739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_157_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10069__I _02330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17467_ _00537_ clknet_leaf_26_clk filters.band\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_172_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14679_ _06669_ _06670_ _06673_ _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__14014__A1 _04728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08492__A2 _00129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16418_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[11\] _08220_ _08225_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14565__A2 _06431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08762__I _01240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17398_ _00468_ clknet_leaf_135_clk channels.env_counter\[1\]\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16349_ _01238_ _01317_ _01334_ channels.exp_counter\[0\]\[4\] _08175_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_89_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15514__A1 channels.sample2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16857__A4 _02847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_1193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_35_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14004__I _05943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13828__A1 _04753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09723_ channels.pw1\[10\] _02091_ _02094_ _02096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09654_ channels.sus_rel3\[6\] _01943_ _01970_ channels.freq1\[14\] _02039_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_179_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08605_ _01113_ _00019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_145_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09585_ channels.atk_dec2\[3\] _01966_ _01972_ _01973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13056__A2 _04905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08536_ _00131_ _01050_ _01036_ _01058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_38_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08467_ net4 _00997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_37_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14005__A1 _04529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09680__A1 channels.atk_dec2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09680__B2 channels.freq3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08672__I _01155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10290__A2 _02385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14556__A2 _06008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_31__f_clk_I clknet_3_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12194__I _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10360_ _01542_ _02541_ _02620_ _02621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_182_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09019_ _01477_ _01478_ _01479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_10291_ _01528_ _02382_ _02549_ _02550_ _02551_ _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_143_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12030_ _04074_ _04090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_72_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09735__A2 _01941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10442__I _02505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13819__A1 _04893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15454__B _07240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13981_ _04631_ _05982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_38_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15720_ _05647_ _07640_ _07333_ _07641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_137_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12932_ _04754_ _04936_ _04937_ _04938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__08847__I _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_124_Left_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15651_ _07574_ _07571_ _07581_ _07583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_107_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12863_ _04868_ _04844_ _04869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_69_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13047__A2 _05049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14244__A1 _04699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14602_ _06515_ _06597_ _06598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11814_ channels.env_counter\[0\]\[8\] channels.env_counter\[1\]\[8\] channels.env_counter\[2\]\[8\]
+ channels.env_counter\[3\]\[8\] _03832_ _01171_ _03905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__15992__A1 _07838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15582_ filters.sample_buff\[5\] _07518_ _07519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12794_ _04443_ _04800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__16285__B _07740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17321_ _00391_ clknet_leaf_87_clk channels.freq1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_28_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14533_ _06455_ _06457_ _06529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_83_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11745_ _03835_ _03836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08474__A2 _01003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_165_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17252_ _00322_ clknet_leaf_18_clk filters.sample_filtered\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_12_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_12_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14464_ _06359_ _06093_ _06461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14547__A2 _05446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11676_ _01168_ _02532_ _03767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16203_ _08057_ _08072_ _08076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12558__A1 _04535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13415_ _05417_ _05420_ _05421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_17183_ _00253_ clknet_leaf_104_clk channels.sus_rel3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10627_ _02835_ _02883_ _02884_ _02885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_36_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09423__A1 _01814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_133_Left_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_14395_ _06189_ _06391_ _06392_ _06393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_141_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08857__S0 _01307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16134_ _07983_ _08008_ _08009_ _07879_ _08010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_141_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09974__A2 _02265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13346_ _04184_ _05351_ _05352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10558_ _02561_ _02776_ _02818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__17547__D _00617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16065_ _07903_ _07914_ _07944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_80_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13277_ _05278_ _05282_ _05283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10489_ _02507_ _02512_ _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15016_ _06962_ _06985_ _06986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12228_ _03255_ _04226_ _04221_ _04234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_121_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_166_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12159_ _03317_ _04164_ _04165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XPHY_EDGE_ROW_142_Left_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_127_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_127_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16967_ _00046_ clknet_leaf_197_clk channels.exp_counter\[1\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15918_ _07785_ _07799_ _07800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_16898_ _00978_ _00844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15027__A3 _06996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15849_ spi_dac_i.counter\[1\] _07720_ spi_dac_i.counter\[2\] _07734_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13038__A2 _04991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09370_ _01770_ _01771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17519_ _00589_ clknet_leaf_22_clk filters.high\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15735__A1 _07650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_151_Left_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_203_clk_I clknet_5_21__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09965__A2 _02265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_218_clk_I clknet_5_21__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14710__A2 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_160_Left_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09706_ _01808_ _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08667__I _01150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_173_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09637_ channels.ctrl_reg2\[5\] _01974_ _01966_ channels.atk_dec2\[5\] _02022_ _02023_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_97_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09568_ filters.cutoff_lut\[11\] _01956_ _01866_ channels.atk_dec3\[2\] _01957_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_65_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08519_ _01041_ _01045_ _01046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_148_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09499_ _01825_ _01853_ _01854_ _01890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09653__A1 filters.cutoff_lut\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11530_ _02328_ _03649_ _03656_ _00405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_18_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_137_Right_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11461_ _03612_ _01515_ _03613_ _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13200_ _05142_ _05147_ _05206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_150_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10412_ _02666_ _02671_ _02672_ _02673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11392_ _03573_ _03569_ _01448_ _03570_ _00350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_14180_ _06176_ _06179_ _06180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_21_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13131_ _05103_ _05109_ _05137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10343_ _02537_ _02545_ _02523_ _02604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_108_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13062_ _03398_ _04219_ _04403_ _05068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_10274_ _02529_ _02532_ _02534_ _02535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_148_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12712__A1 _04701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12013_ _04010_ _04076_ _04080_ _00464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_1193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_109_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16821_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[2\] _00916_ _00920_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_144_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14465__A1 _05509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16752_ _03710_ _00868_ _00870_ _00806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11279__A1 filters.cutoff_lut\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13964_ _05762_ _05964_ _05965_ _05966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_161_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15703_ _07626_ _00608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12915_ _04918_ _04919_ _04920_ _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_16683_ _08421_ _08424_ _08281_ _08426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_17_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13895_ _05890_ _05896_ _05897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_115_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15634_ channels.sample1\[9\] _03427_ _07567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12846_ _04733_ _04849_ _04851_ _04852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_75_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_158_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15565_ channels.sample1\[4\] _03400_ _07503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_167_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12777_ filters.cutoff_lut\[12\] _04442_ _04783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09644__A1 filters.res_filt\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09644__B2 _02029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17304_ _00374_ clknet_leaf_152_clk channels.accum\[1\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14516_ _06304_ _06395_ _06494_ _06511_ _06512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_11728_ _03817_ _03818_ _03757_ _03819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15496_ filters.low\[31\] _07428_ _07439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_182_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17235_ _00305_ clknet_leaf_171_clk channels.sample1\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14447_ _06438_ _06443_ _06444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_104_Right_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11659_ _03747_ _03749_ _03750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_17166_ _00236_ clknet_leaf_143_clk channels.ctrl_reg3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14378_ _06374_ _06375_ _06376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14940__A2 _06912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_101_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_168_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16117_ _07991_ _07993_ _07994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12951__A1 _04456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13329_ _05333_ _05254_ _05334_ _05335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_49_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17097_ _00167_ clknet_leaf_99_clk channels.ctrl_reg1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_10_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_1_0_clk clknet_0_clk clknet_3_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_16048_ _07760_ _07875_ _07927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_0_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_161_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09255__S0 _01144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12703__A1 _04265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08870_ _01339_ _01340_ _01341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_122_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_181_3738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_3749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14456__A1 _06337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09422_ filters.hp _01803_ _01809_ _01815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11690__A1 channels.sus_rel3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15956__A1 _07598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11690__B2 channels.sus_rel2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_99_clk_I clknet_5_13__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09353_ net9 _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_19_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_142_clk_I clknet_5_30__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10245__A2 _02505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09284_ channels.lfsr\[0\]\[20\] _01712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_22_clk_I clknet_5_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10257__I _01141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_157_clk_I clknet_5_29__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14931__A2 _04160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_37_clk_I clknet_5_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16684__A2 _08244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09246__S0 _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14695__A1 _03411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_89_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08999_ _01460_ _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_138_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_3_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09323__B1 _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16828__B _01823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_67_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10961_ _03185_ _03186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09874__A1 channels.ctrl_reg2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13670__A2 _05671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12700_ _04705_ _04268_ _04706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_168_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13680_ _04512_ _04447_ _05481_ _05684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_57_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_84_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10892_ _02056_ _03105_ _03142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_167_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12631_ _03256_ _04566_ _04633_ _04634_ _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_155_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_100_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09626__A1 channels.freq1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09626__B2 channels.pw3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13422__A2 _05415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10236__A2 channels.ctrl_reg3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15350_ _07303_ _07304_ _07305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_81_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12562_ _04565_ _04567_ _04568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_80_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16563__B _08292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14301_ _06168_ _06278_ _06299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11513_ channels.pw1\[1\] _03643_ _03644_ _03646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_124_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_108_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15281_ _07235_ _07239_ _07241_ _07242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_136_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12493_ _04292_ _04498_ _04423_ _04499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_110_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17020_ _00099_ clknet_leaf_232_clk channels.lfsr\[2\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_22_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14232_ _06150_ _06155_ _06231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11444_ _01219_ _03604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12933__A1 _04846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14163_ _06085_ _06162_ _06163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_61_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11375_ channels.accum\[2\]\[4\] _03563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_150_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13114_ _04888_ _04889_ _05120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_104_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10326_ _01598_ _02385_ _02587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14094_ _05446_ _06093_ _06010_ _06094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09237__S0 _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13045_ _04928_ _04930_ _05051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_163_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10257_ _01141_ _02518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10188_ channels.pw1\[5\] _02435_ _02449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16804_ _01741_ _00906_ _00908_ _00901_ _00820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_17784_ _00854_ clknet_leaf_215_clk channels.exp_periods\[0\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14996_ _06961_ _06966_ _06967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_89_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13110__A1 _04902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16735_ _03710_ _08464_ _08466_ _00800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_117_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13947_ _04238_ _04847_ _05279_ _05947_ _05949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_89_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09865__A1 channels.ctrl_reg2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16666_ _08406_ _08410_ _08292_ _08412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11672__A1 channels.sus_rel3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11672__B2 channels.sus_rel2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13878_ _05785_ _05844_ _05880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_72_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15617_ _03372_ _07549_ _07550_ _03395_ _07551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_147_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12829_ _04316_ _04480_ _04835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16597_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[9\] _08370_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[9\]
+ _08371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15548_ filters.sample_buff\[2\] _07478_ _07487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_29_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14772__I _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15479_ _07422_ _07423_ _00587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_150_clk clknet_5_29__leaf_clk clknet_leaf_150_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_16_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15166__A2 channels.sample1\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17218_ _00288_ clknet_leaf_174_clk channels.sample2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12924__A1 _04295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17149_ _00219_ clknet_leaf_142_clk channels.sus_rel2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_141_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09971_ _02098_ _02266_ _02271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08922_ _01387_ _01388_ _01389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_0_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09553__B1 _01941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08853_ channels.freq3\[1\] _01074_ _01325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14429__A1 _05721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11636__I _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08784_ _01257_ _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_97_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16648__B _08313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09856__A1 _02098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11663__A1 _03535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09405_ _01017_ _01800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_45_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09608__A1 channels.ctrl_reg2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09608__B2 channels.atk_dec2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09336_ net8 _01739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_164_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_168_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15778__I _07630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09267_ _01626_ _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_141_clk clknet_5_30__leaf_clk clknet_leaf_141_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_161_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08680__I _01163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09198_ channels.lfsr\[2\]\[8\] _01639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_105_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11160_ _03375_ _03376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14668__A1 _06456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_8_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10111_ _02371_ _02372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_179_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11091_ _03189_ _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_140_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10042_ _02309_ _02321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13340__A1 _05341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11546__I _02149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10450__I _02505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14850_ _06797_ _06831_ _06832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_26_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13801_ _04705_ _05260_ _05804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14781_ _06769_ _06756_ _06770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11993_ _04044_ _04063_ _04064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16520_ _08274_ _08305_ _08306_ _08307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_97_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13732_ _05728_ _05735_ _05736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_86_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10944_ _03168_ _03080_ _03173_ _00302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_129_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16451_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[3\] _08247_ _08098_ _08250_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13663_ _05584_ _05600_ _05667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__16593__A1 _08238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10875_ _03118_ _03116_ _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_168_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_156_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15402_ _07351_ _07352_ _07353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_27_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12614_ _04615_ _04619_ _04620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16382_ _08197_ _08198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13594_ _05594_ _05598_ _05599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_66_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09075__A2 _01334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_156_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15333_ _07288_ _07289_ _00575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_109_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12545_ _04549_ _04547_ _04550_ _04551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
Xclkbuf_leaf_132_clk clknet_5_31__leaf_clk clknet_leaf_132_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_137_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13159__A1 _05138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15264_ _05751_ _07219_ _07217_ _07225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_123_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12476_ _04478_ _04479_ _04481_ _04482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_0_151_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12906__A1 _04833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17003_ _00082_ clknet_leaf_218_clk channels.lfsr\[2\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14215_ _06211_ _06212_ _06213_ _06214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_22_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_5 _01590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11427_ channels.accum\[1\]\[1\] _03593_ _03594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15195_ _01747_ channels.sample1\[9\] _07159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_134_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14146_ _06144_ _06145_ _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_1_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11358_ _01254_ _03551_ _01931_ _03552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_162_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10309_ channels.ch3_env\[6\] _02570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_130_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14077_ _06072_ _06077_ _06078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__15320__A2 _06065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11289_ net15 _03494_ _03495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_67_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13331__A1 _05234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13028_ _04435_ _04518_ _05033_ _05034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11893__A1 _03128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer17 _06063_ net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09838__A1 channels.freq2\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrebuffer28 _04235_ net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_17767_ _00837_ clknet_leaf_201_clk channels.exp_periods\[2\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_178_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer39 _04388_ net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_88_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14979_ _06935_ _06950_ _06951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_107_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16718_ _08445_ _08454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17698_ _00768_ clknet_leaf_222_clk channels.lfsr\[0\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_176_3648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_176_3659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16584__A1 _08356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16649_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[1\] _08397_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_147_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13398__A1 _05403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09121_ _01300_ _01570_ _01571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_123_clk clknet_5_30__leaf_clk clknet_leaf_123_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_5_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16336__A1 _03974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09052_ _01509_ _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_114_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14898__A1 _06614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12373__A2 _04378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09954_ channels.freq3\[13\] _02258_ _02255_ _02260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15311__A2 _06910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13322__A1 _04315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08905_ _01367_ _01368_ _01373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09885_ channels.atk_dec2\[0\] _02211_ _02206_ _02212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12676__A3 _04675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13873__A2 _05848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08836_ _01308_ channels.accum\[1\]\[0\] _01309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15282__B _06899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08767_ channels.exp_counter\[2\]\[2\] _01090_ _01228_ _01241_ _01244_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09829__A1 channels.freq2\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13625__A2 _04884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08698_ _01179_ _01180_ _01181_ _01173_ _01182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_178_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_24_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10660_ _02662_ _02872_ _02918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09319_ _01663_ _01732_ _01733_ _01666_ _00113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_114_clk clknet_5_26__leaf_clk clknet_leaf_114_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_146_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10591_ _02848_ _02807_ _02849_ _02850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_63_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12330_ _03287_ _04219_ _04196_ _04336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_17_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_151_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12261_ _03348_ _04190_ _04267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_TAPCELL_ROW_151_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14000_ _05950_ _05954_ _06001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__12364__A2 _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11212_ _03423_ _03424_ _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput20 net20 DAC_dat_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_12192_ filters.res_lut\[4\] _04168_ _04198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_TAPCELL_ROW_112_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11143_ filters.low\[8\] _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_112_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15951_ _07764_ _07832_ _07833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10127__A1 _01534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11074_ _03293_ _03295_ _03296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11276__I _02334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10025_ _02104_ _02308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14902_ _06851_ _06879_ _06880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_15882_ _07747_ _07753_ _07763_ _07764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15066__A1 _07032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08740__A1 _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17621_ _00691_ clknet_leaf_128_clk channels.env_counter\[3\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14833_ _06795_ _06800_ _06808_ _06816_ _06817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_53_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11627__A1 channels.pw2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08585__I _01100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14764_ _06700_ _06754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_17552_ _00622_ clknet_leaf_14_clk filters.low\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11976_ _03843_ _04045_ _04050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_158_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_158_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16503_ _08285_ _08290_ _08292_ _08293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13715_ _05623_ _05634_ _05718_ _05719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_17483_ _00553_ clknet_leaf_244_clk filters.band\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10927_ _03162_ _02783_ _03163_ _00295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14695_ _03411_ _03221_ _06690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16434_ tt_um_rejunity_sn76489.clk_counter\[2\] tt_um_rejunity_sn76489.clk_counter\[1\]
+ tt_um_rejunity_sn76489.clk_counter\[0\] _08236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_13646_ _05548_ _05650_ _05651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_160_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10858_ _03089_ _03090_ _03110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__14041__A2 _06041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16365_ channels.ch3_env\[4\] _08185_ _08186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_105_clk clknet_5_15__leaf_clk clknet_leaf_105_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_26_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13577_ _05508_ _05521_ _05581_ _05582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_87_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10789_ _03021_ _03022_ _03043_ _03044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_171_3556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15316_ _07246_ _07249_ _07274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_17__f_clk clknet_3_4_0_clk clknet_5_17__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10602__A2 _02622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12528_ _04172_ _04210_ _04534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_16296_ _08145_ _00682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_136_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_132_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15247_ _07184_ _07185_ _07209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_132_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12459_ _04463_ _04408_ _04464_ _04465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_22_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_8__f_clk_I clknet_3_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15178_ _07139_ _07141_ _07142_ _07143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14129_ _04376_ _05077_ _06129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10118__A1 _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09670_ _02042_ _02053_ _02054_ _00147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_118_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_19_Left_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08621_ _01121_ _00027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13607__A2 _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08552_ _01062_ _01068_ _01069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__11618__A1 _03664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16926__B _00877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16557__A1 _08333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08483_ _01004_ _01013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_76_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12745__I _04750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_28_Left_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09104_ _01555_ _01556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_94_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08798__A1 channels.ctrl_reg3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13791__A1 _04525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09035_ _01492_ _01493_ _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_96_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15532__A2 _07468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12897__A3 _04450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09937_ _02246_ _02248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_102_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_37_Left_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13846__A2 _05848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09868_ channels.ctrl_reg2\[3\] _02195_ _02199_ _02200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_70_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08819_ _01291_ _01292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09799_ _02149_ _02150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_29_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11830_ _03915_ _03920_ _03921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11609__A1 _01780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16836__B _00877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11761_ _03837_ _03839_ _03824_ _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13500_ _04401_ _05505_ _05506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10712_ _02949_ _02951_ _02968_ _02969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_95_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14480_ _06353_ _06368_ _06477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11692_ _01277_ _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_126_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13431_ _05374_ _05437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_153_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10643_ _02590_ _02637_ _02901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_153_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16150_ _08010_ _08025_ _08026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_153_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13362_ _04596_ _05367_ _05262_ _05368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_106_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10574_ _02830_ _02833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_107_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__16571__B _08301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer8 _05031_ net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15101_ _07040_ _07050_ _07068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_114_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12313_ _04313_ _04318_ _04319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_77_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16081_ _07930_ _07881_ _07804_ _07959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_107_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16720__A1 _08453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13293_ _05296_ _05297_ _05298_ _05299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_45_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15032_ _06971_ _06974_ _07002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_107_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12244_ _04234_ _04239_ _04250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12390__I _04395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12175_ _04180_ _04181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_11126_ _03228_ _03344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_16983_ _00062_ clknet_leaf_168_clk channels.accum\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15934_ _07813_ _07814_ _07815_ _07816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_11057_ _03278_ _03279_ _03280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15039__A1 _05969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10008_ channels.atk_dec3\[2\] _02292_ _02294_ _02297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15865_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[3\] _07746_ _07747_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_161_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17604_ _00674_ clknet_leaf_44_clk net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_14816_ _06748_ _06801_ _06802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_125_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15796_ filters.low\[22\] _07694_ _07695_ _07696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_157_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17535_ _00605_ clknet_leaf_200_clk channels.exp_periods\[3\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11959_ _03854_ _04032_ _04036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_114_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14747_ _03456_ _06508_ _06738_ _06610_ _00540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_114_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14678_ _06671_ _06672_ _06673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17466_ _00536_ clknet_5_1__leaf_clk filters.band\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15211__A1 _03394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_55_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16417_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[10\] _08223_ _08224_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_157_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13629_ _05629_ _05633_ _05634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_17397_ _00467_ clknet_leaf_131_clk channels.env_counter\[1\]\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13773__A1 _04597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16348_ _08174_ _00705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16279_ _08136_ _08137_ _00673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_164_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16711__A1 _03710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13525__A1 _05527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12879__A3 _04884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09722_ _01757_ _02090_ _02095_ _00158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_52_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09653_ filters.cutoff_lut\[15\] _01988_ _02038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10511__A1 _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08604_ channels.lfsr\[3\]\[6\] _01113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_179_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09584_ _01967_ _01968_ _01969_ _01971_ _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_145_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_118_Right_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_179_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08535_ _01030_ _00131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12264__A1 _04266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13764__A1 _04667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09018_ channels.freq2\[13\] _01279_ _01293_ channels.freq1\[13\] _01478_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__13516__A1 _05508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10290_ _01615_ _02385_ _02551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_176_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13980_ _05560_ _05980_ _05894_ _05981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_146_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12931_ _04644_ _04759_ _04757_ _04937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_88_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15650_ _07574_ _07571_ _07581_ _07582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_12862_ _04867_ _04846_ _04868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_107_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15441__A1 _07373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16566__B _08339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11813_ _03902_ _03903_ _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14601_ _06517_ _06596_ _06597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_96_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12255__A1 _03288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15581_ _07516_ _07517_ _07518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_179_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12793_ _04787_ _04798_ _04799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09120__A1 _01086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17320_ _00390_ clknet_leaf_77_clk channels.freq1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14532_ _06455_ _06457_ _06528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11744_ _03823_ _03835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_84_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17251_ _00321_ clknet_leaf_86_clk filters.sample_filtered\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14463_ _06363_ _06364_ _06459_ _06460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_166_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11675_ channels.sus_rel2\[7\] _01281_ _01295_ channels.sus_rel1\[7\] _03765_ _03766_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_12_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_12_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16202_ _08074_ _08075_ _00658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13414_ _04775_ _05418_ _05419_ _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__12558__A2 _04537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17182_ _00252_ clknet_leaf_106_clk channels.sus_rel3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10626_ _02837_ _02878_ _02884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_70_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14394_ _06192_ _06274_ _06392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_84_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08857__S1 _01328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16133_ _07757_ _07955_ _08009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13345_ _05350_ _05351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_134_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10557_ _02755_ _02760_ _02758_ _02817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_52_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13507__A1 _05512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16064_ _07929_ _07938_ _07942_ _07943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_13276_ _04302_ _05281_ _05282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10488_ _02592_ _02528_ _02576_ _02749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_15015_ _06964_ _06965_ _06985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12227_ _04223_ _04232_ _04233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_121_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_166_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12158_ _04163_ _04164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_11109_ _03242_ _03328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12089_ _04064_ _04104_ _04125_ _00495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16966_ _00045_ clknet_leaf_196_clk channels.exp_counter\[1\]\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_127_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14483__A2 _05563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15917_ _07797_ _07798_ _07799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16897_ _00966_ channels.exp_periods\[1\]\[2\] _00975_ _00978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11464__I _01219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15848_ spi_dac_i.counter\[2\] spi_dac_i.counter\[1\] _07720_ _07733_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_152_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15432__A1 _06934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15779_ _03733_ _07683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17518_ _00588_ clknet_leaf_37_clk filters.high\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_157_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_144_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12295__I _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17449_ _00519_ clknet_leaf_190_clk channels.accum\[3\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_156_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_101_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10980__A1 _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11639__I _01750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_54_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15671__A1 _03239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09705_ _01801_ _02081_ _02083_ _00153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11288__A2 _01093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_94_clk clknet_5_7__leaf_clk clknet_leaf_94_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09636_ _01908_ _02019_ _02020_ _02021_ _02022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_97_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_179_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09567_ _01851_ _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_139_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08518_ _01024_ _01027_ _01044_ _01045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__08683__I _01166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09498_ _01875_ _01878_ _01883_ _01888_ _01889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_33_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10718__I _02974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11460__A2 _03605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16833__C _04101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11460_ channels.accum\[1\]\[15\] _03605_ _03613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10411_ _02669_ _02670_ _02672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11391_ channels.accum\[2\]\[10\] _03573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13130_ _05113_ _05136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10342_ _02599_ _02600_ _02602_ _02603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_131_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13061_ _04705_ _04751_ _05067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10273_ _01156_ _02533_ _02534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_148_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12012_ channels.env_counter\[1\]\[0\] _04079_ _04080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_148_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16820_ _01756_ _00915_ _00918_ _00919_ _00825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__17162__CLK clknet_5_26__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_109_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15662__A1 filters.sample_buff\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16751_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[4\] _00869_ _00863_ _00870_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13963_ _05765_ _05845_ _05965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11284__I net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_161_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_85_clk clknet_5_12__leaf_clk clknet_leaf_85_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15702_ channels.exp_periods\[3\]\[3\] _07626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12914_ _04237_ _04273_ _04920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16682_ _08421_ _08424_ _08425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13894_ _05894_ _05895_ _05896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_17_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12845_ _04848_ _04850_ _04268_ _04181_ _04851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_15633_ channels.sample2\[9\] _03424_ _07565_ _03233_ _07566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_29_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12776_ _03200_ _04216_ _04781_ _04782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_61_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15564_ channels.sample2\[4\] _03377_ _07501_ _03230_ _07502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_127_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17303_ _00373_ clknet_leaf_163_clk channels.accum\[1\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11727_ channels.sus_rel3\[3\] _03782_ _03783_ channels.sus_rel2\[3\] _03818_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_139_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14515_ _06495_ _06509_ _06510_ _06511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_138_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15495_ _07430_ _07437_ _07438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__11451__A2 _03605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17234_ _00304_ clknet_leaf_171_clk channels.sample1\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14446_ _06439_ _06442_ _06443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_11658_ _03748_ _03742_ _03749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_37_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10609_ _02866_ _02867_ _02868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_17165_ _00235_ clknet_leaf_144_clk channels.ctrl_reg3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14377_ _06233_ _06250_ _06375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11834__S0 _03886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11589_ channels.pw3\[0\] _03697_ _03698_ _03699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16116_ _07776_ _07992_ _07993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_168_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13328_ _05255_ _05263_ _05334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17096_ _00166_ clknet_leaf_99_clk channels.ctrl_reg1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11459__I _02364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16047_ _07916_ _07918_ _07925_ _07926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13259_ _05244_ _05247_ _05264_ _05265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_86_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09255__S1 _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13900__A1 _05813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_181_3739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09580__A1 filters.mode_vol\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09580__B2 channels.sus_rel2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15653__A1 filters.sample_buff\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16949_ _00028_ clknet_leaf_238_clk channels.lfsr\[3\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_76_clk clknet_5_14__leaf_clk clknet_leaf_76_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09332__A1 _01710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09421_ _01813_ _01814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_17_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12482__A4 _03410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09352_ _01742_ _01743_ _01754_ _00125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_19_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_47_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12234__A4 filters.high\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09283_ channels.lfsr\[2\]\[21\] _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_157_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13719__A1 _03398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13195__A2 _05157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14392__A1 _06305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12753__I _04758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16225__I _07683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14144__A1 _04742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09246__S1 _01680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14695__A2 _03221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09571__A1 channels.freq1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09571__B2 channels.freq3\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08678__I _01161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_10_Left_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08998_ _01256_ _01460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_138_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10181__A2 _01286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_67_clk clknet_5_11__leaf_clk clknet_leaf_67_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_138_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_170_Right_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10960_ _03184_ _03185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_104_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09619_ _01998_ _02000_ _02002_ _02005_ _02006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_10891_ _03125_ _03135_ _03139_ _03140_ _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_167_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12630_ _04615_ _04632_ _04635_ _04636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_38_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16844__B _00877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12561_ _03255_ _04566_ _04504_ _04567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_65_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11512_ _03639_ _03642_ _03645_ _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14300_ _06295_ _06296_ _06297_ _06183_ _06298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_80_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15280_ _07235_ _07239_ _07240_ _07241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_163_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12492_ _04416_ _04498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_164_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14231_ _06197_ _06229_ _06230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_22_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11443_ _01104_ _03603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_135_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17528__CLK clknet_5_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14162_ _06101_ _06161_ _06162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_11374_ _03138_ _01359_ _03562_ _00343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13113_ _04888_ _04889_ _05119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10325_ _01510_ _02377_ _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_14093_ _06005_ _06093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09972__I _02101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09237__S1 _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13044_ _04928_ _04930_ _05050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10256_ _01306_ channels.env_vol\[3\]\[2\] _02516_ _02517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_163_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_163_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09562__A1 channels.ctrl_reg2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09562__B2 channels.freq2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10187_ _01265_ _01263_ channels.pw2\[5\] _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_56_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16803_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[0\] _00907_ _00908_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_202_clk_I clknet_5_21__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17783_ _00853_ clknet_leaf_214_clk channels.exp_periods\[0\]\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_58_clk clknet_5_8__leaf_clk clknet_leaf_58_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_14995_ _06964_ _06965_ _06966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_156_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13110__A2 _04903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16734_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[4\] _08465_ _08459_ _08466_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13946_ _04238_ _05279_ _05947_ _04847_ _05948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_159_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16665_ _08406_ _08410_ _08411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13877_ _05769_ _05781_ _05878_ _05879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_159_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_217_clk_I clknet_5_21__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13949__A1 _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15616_ channels.sample3\[8\] _07538_ _07550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12828_ _04324_ _04729_ _04834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_16596_ _08242_ _08329_ _08370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_178_3690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15547_ _07449_ _07486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_139_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12759_ _04764_ _04765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15478_ filters.high\[29\] _06983_ _07333_ _07423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17217_ _00287_ clknet_leaf_174_clk channels.sample2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14429_ _05721_ _05079_ _06426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_170_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11807__S0 _01150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12924__A2 _04929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17148_ _00218_ clknet_leaf_145_clk channels.sus_rel2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_40_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09970_ channels.pw3\[11\] _02270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_110_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17079_ _00149_ clknet_leaf_107_clk channels.freq1\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08921_ channels.freq2\[6\] _01276_ _01289_ channels.freq1\[6\] _01388_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09553__A1 channels.pw1\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09553__B2 channels.ctrl_reg1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08852_ _01160_ _01310_ _01313_ _01303_ _01324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_100_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08783_ _01256_ _01257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_49_clk clknet_5_10__leaf_clk clknet_leaf_49_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09305__A1 _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09404_ _01777_ _01793_ _01799_ _00136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_95_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09069__B1 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09335_ _01720_ _01722_ _01726_ _01738_ _00124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10268__I _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09266_ _01695_ _01696_ _01690_ _01697_ _01679_ _01680_ _01698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_118_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13168__A2 _04737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14365__A1 _05509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09197_ _01633_ _01634_ _01638_ _01627_ _00086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_62_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10926__A1 channels.sample1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15794__I _07630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14117__A1 _04803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09792__A1 _02110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10110_ _01264_ _02369_ _02370_ _02371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11090_ filters.low\[5\] _03310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10041_ _02309_ _02320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13340__A2 _05345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11351__A1 _01585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13800_ _05697_ _05801_ _05802_ _05803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_98_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11992_ _03911_ _04059_ _04063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_14780_ _06768_ _06769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13731_ _05729_ _05734_ _05735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10943_ channels.sample1\[7\] _03170_ _03173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12851__A1 _04853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16450_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[3\] _08247_ _08249_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13662_ _05664_ _05665_ _05666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10874_ _03109_ _03120_ _03124_ _03125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xclkbuf_3_0_0_clk clknet_0_clk clknet_3_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_27_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15401_ filters.low\[23\] _06701_ _07352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_112_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12613_ _04498_ _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10178__I channels.pw1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16381_ tt_um_rejunity_sn76489.noise\[0\].gen.signal_edge.previous_signal_state_0
+ _02349_ _08197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_13593_ _05595_ _05596_ _05597_ _05598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_26_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_156_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12544_ _04545_ _04546_ _04550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15332_ filters.high\[17\] _07033_ _06899_ _07289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_137_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16345__A2 _01317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10090__A1 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13489__I _05341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14356__A1 filters.band\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12475_ _04220_ _04480_ _04481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15263_ _07035_ _07222_ _07224_ _00570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_117_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17002_ _00081_ clknet_leaf_218_clk channels.lfsr\[2\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_152_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12906__A2 _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14214_ _04896_ _05181_ _06213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_11426_ _03149_ _03593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_6 _01590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09232__B1 _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15194_ _01761_ channels.sample2\[9\] _07158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_134_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09783__A1 _01814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14145_ filters.band\[26\] _04186_ _06145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11357_ _03546_ _03549_ _03550_ _03551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__11590__A1 _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10308_ _02567_ _02538_ _02568_ _02569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_67_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_98_clk_I clknet_5_13__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14076_ _06074_ _06076_ _06077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11288_ _01824_ _01093_ _01831_ _03493_ _03494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_13027_ _04438_ _04517_ _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_clkbuf_leaf_141_clk_I clknet_5_30__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09535__B2 channels.pw3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10239_ _02372_ _02379_ _02388_ _02499_ _02500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_20_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_21_clk_I clknet_5_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11673__S _03763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09651__B _02036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17766_ _00836_ clknet_leaf_58_clk tt_um_rejunity_sn76489.clk_counter\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xrebuffer18 _05330_ net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer29 _04880_ net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14978_ _06938_ _06949_ _06950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA_clkbuf_leaf_156_clk_I clknet_5_29__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16717_ _01765_ _08453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11645__A2 _03728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10448__A3 _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13929_ _05828_ _05930_ _05931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17697_ _00767_ clknet_leaf_221_clk channels.lfsr\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16648_ _08395_ _08396_ _08313_ _00783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_176_3649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13398__A2 _05379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16579_ _08135_ _08356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_123_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_174_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09120_ _01086_ _01569_ _01570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08781__I _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09051_ _01508_ _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_170_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_142_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10908__A1 channels.sample2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15847__A1 _07598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09953_ _02234_ _02257_ _02259_ _00225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_109_clk_I clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09526__A1 _01913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08904_ _01362_ _01262_ _01372_ _01318_ _00059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_110_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09884_ _02209_ _02211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08835_ _01307_ _01308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__16272__A1 filters.sample_buff\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08766_ _01243_ _00050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08956__I _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input11_I bus_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_25__f_clk_I clknet_3_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08697_ _01176_ channels.exp_periods\[3\]\[0\] _01181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15789__I _07663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09318_ _01657_ _01732_ _01733_ _01661_ _00112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_180_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08691__I _01152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10590_ _02713_ _02750_ _02805_ _02847_ _02849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_91_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10072__A1 filters.cutoff_lut\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14338__A1 _06211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11331__B _03517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09249_ _01610_ _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_181_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12260_ _04265_ _04266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_79_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13010__A1 _04993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_151_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_151_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11211_ _03395_ _03424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11021__B1 _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12191_ _04196_ _04197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_181_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput21 net21 DAC_le vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__11572__A1 _03666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11142_ filters.high\[8\] _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_112_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14510__A1 _06403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15950_ _07807_ _07831_ _07832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11073_ _03294_ _03278_ _03295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_179_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10024_ _02242_ _02301_ _02307_ _00248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14901_ _06874_ _06878_ _06879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_15881_ _07762_ _07763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_17620_ _00690_ clknet_leaf_147_clk channels.env_counter\[3\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14832_ _06794_ _06807_ _06765_ _06816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_153_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13616__A3 _04804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17551_ _00621_ clknet_leaf_14_clk filters.low\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14763_ _06752_ _06753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_11975_ _04043_ _04047_ _04049_ _00457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16502_ _08257_ _08292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_158_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_158_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13714_ _05629_ _05633_ _05718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17482_ _00552_ clknet_leaf_244_clk filters.band\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10926_ channels.sample1\[0\] _01560_ _03163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14694_ _06688_ _06689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_85_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09128__S0 _01201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16433_ tt_um_rejunity_sn76489.clk_counter\[4\] tt_um_rejunity_sn76489.clk_counter\[3\]
+ _08235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10857_ _03099_ _03101_ _03109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13645_ _05646_ _05649_ _05650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_67_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16364_ _08178_ _08185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_136_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13576_ _05580_ _05520_ _05581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10788_ _03025_ _03042_ _03043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_137_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_171_3557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10063__A1 filters.cutoff_lut\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14329__A1 _04806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15315_ _07271_ _07254_ _07263_ _07264_ _07273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_26_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12527_ _04532_ _04528_ _04533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16295_ channels.env_counter\[3\]\[3\] _08145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_87_1164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_132_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15246_ _07184_ _07185_ _07208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12458_ _04383_ _04394_ _04464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_140_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09756__A1 channels.ctrl_reg1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11409_ _03583_ _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_111_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12389_ _03381_ _04341_ _04395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_15177_ _07139_ _07141_ _07086_ _07142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15829__A1 _07598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14128_ _06037_ _06126_ _06127_ _06128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10371__I channels.ch3_env\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14059_ _05882_ _05961_ _06060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11315__A1 _03513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input3_I addr[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_68_Right_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_158_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08620_ channels.lfsr\[3\]\[14\] _01121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_178_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08551_ clk_trg\[1\] _01064_ _01067_ clk_trg\[0\] _01068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_89_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17749_ _00819_ clknet_leaf_55_clk tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08482_ net14 _01011_ _01012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_76_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14568__A1 _04355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_77_Right_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13240__A1 _05157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09103_ channels.accum\[0\]\[21\] channels.accum\[1\]\[21\] channels.accum\[2\]\[21\]
+ channels.accum\[3\]\[21\] _01139_ _01480_ _01555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__10054__A1 _02328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09995__A1 _02240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09034_ channels.freq2\[14\] _01280_ _01293_ channels.freq1\[14\] _01493_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_131_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_96_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_96_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09747__A1 channels.ctrl_reg1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14740__A1 _06703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11554__A1 _03673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_86_Right_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13793__S _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08970__A2 _01360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09936_ _02246_ _02247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10109__A2 channels.ctrl_reg3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09867_ _02175_ _02199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_70_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16245__A1 _07923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08818_ _01290_ _01291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08686__I _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13059__A1 _04699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09798_ _01017_ _02149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_73_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_29_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08749_ _01103_ _01230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_5_23__f_clk clknet_3_5_0_clk clknet_5_23__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_95_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11760_ _03837_ _03850_ _03851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_166_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16548__A2 _08267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10711_ _02959_ _02967_ _02968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_95_Right_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_113_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11691_ _01397_ _03782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15220__A2 channels.sample3\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13430_ _05299_ _05358_ _05436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10642_ _02501_ _02601_ _02900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_153_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_180_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10045__A1 _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09986__A1 _02215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13361_ _05187_ _05367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_107_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10573_ _02359_ _02831_ _02832_ _00272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15100_ _07043_ _07049_ _07067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12312_ _04317_ _04318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xrebuffer9 net37 net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16080_ _07811_ _07829_ _07957_ _07958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_13292_ _05203_ _05241_ _05298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15468__B _07356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09738__A1 channels.ctrl_reg1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12243_ _04246_ _04247_ _04248_ _04249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_15031_ _06997_ _07000_ _07001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_20_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12337__A3 _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11545__A1 _03666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12888__A4 _04378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12174_ _04179_ _04180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_2_Left_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11125_ filters.high\[7\] _03343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_120_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13298__A1 _05211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16982_ _00061_ clknet_leaf_188_clk channels.accum\[0\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15933_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[0\] _07812_ _07815_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11056_ _03267_ _03261_ _03277_ _03279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_155_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09910__A1 channels.sus_rel2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10007_ _02250_ _02291_ _02296_ _00242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_129_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15864_ _07745_ _07746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_17603_ _00673_ clknet_leaf_41_clk spi_dac_i.spi_dat_buff_0\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14798__A1 filters.band\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14815_ _06795_ _06800_ _06801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_15795_ _07683_ _07695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_125_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17534_ _00604_ clknet_leaf_20_clk filters.sample_buff\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14746_ _06403_ _06737_ _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08477__A1 _01006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11958_ _04027_ _04034_ _04035_ _00454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17465_ _00535_ clknet_leaf_2_clk filters.band\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10909_ _03147_ _03013_ _03152_ _00288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14677_ _06580_ _06588_ _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11889_ channels.env_vol\[0\]\[5\] _03965_ _03975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15211__A2 _07162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16416_ _08190_ _08223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_15_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13628_ _05630_ _05631_ _05632_ _05633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_55_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17396_ _00466_ clknet_leaf_132_clk channels.env_counter\[1\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10036__A1 channels.sus_rel3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16347_ _01235_ _01317_ _01334_ channels.exp_counter\[0\]\[3\] _08174_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_13559_ _05563_ _05370_ _05453_ _05564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_42_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16278_ filters.sample_buff\[14\] _07742_ _08116_ spi_dac_i.spi_dat_buff_0\[10\]
+ spi_dac_i.spi_dat_buff_0\[11\] _08096_ _08137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_140_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_164_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13525__A2 _05530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15229_ _07176_ _07191_ _07192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__11536__A1 _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09721_ channels.pw1\[9\] _02091_ _02094_ _02095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_52_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11839__A2 _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09901__A1 _02155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09652_ _02023_ _02035_ _02037_ _00146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_59_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08603_ _01112_ _00018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_171_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09583_ channels.pw3\[11\] _01841_ _01970_ channels.freq1\[11\] _01971_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15450__A2 _06734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08534_ _01021_ _01055_ _01056_ _01057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_77_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_171_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13461__A1 _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12264__A2 _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09968__A1 channels.pw3\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16702__A2 _08437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09017_ channels.freq3\[13\] _01079_ _01477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14713__A1 _06706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11527__A1 channels.pw1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_72_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09919_ _02149_ _02234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_146_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12930_ _04632_ _04759_ _04757_ _04936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_69_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12861_ _04852_ _04857_ _04866_ _04867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_77_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_107_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14600_ _06519_ _06595_ _06596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_11812_ channels.env_counter\[0\]\[7\] channels.env_counter\[1\]\[7\] channels.env_counter\[2\]\[7\]
+ channels.env_counter\[3\]\[7\] _01151_ _03842_ _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_15580_ channels.sample1\[5\] _03401_ _07517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12792_ _04790_ _04797_ _04798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_69_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14531_ _06484_ _04631_ _06527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11743_ _03830_ _03833_ _03834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_166_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17250_ _00320_ clknet_5_6__leaf_clk filters.sample_filtered\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14462_ _04576_ _05990_ _06365_ _06459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11674_ channels.sus_rel3\[7\] _01080_ _03765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_126_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_12_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16582__B _08301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10018__A1 _02234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16201_ spi_dac_i.spi_dat_buff_1\[7\] _07719_ _07870_ spi_dac_i.spi_dat_buff_1\[8\]
+ _07871_ _08075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_37_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13413_ _04874_ _04951_ _05419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_17181_ _00251_ clknet_leaf_72_clk channels.sus_rel3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10625_ _02879_ _02883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14393_ _06192_ _06274_ _06391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16132_ _07757_ _07955_ _07843_ _08008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10556_ _02797_ _02815_ _02816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13344_ filters.high\[19\] filters.band\[19\] _04710_ _05350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_84_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13507__A2 _05510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16063_ _07825_ _07823_ _07939_ _07940_ _07941_ _07942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_13275_ _05280_ _05281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10487_ _02592_ _02543_ _02638_ _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_51_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11518__A1 _03515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15014_ _06944_ _06946_ _06967_ _06966_ _06961_ _06984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_122_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12226_ _03255_ _04226_ _04231_ _04232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__14180__A2 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_244_clk clknet_5_0__leaf_clk clknet_leaf_244_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_166_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12157_ _04162_ _04163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_166_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11108_ _03244_ _03327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12088_ channels.env_counter\[0\]\[12\] _04107_ _04125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_159_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16965_ _00044_ clknet_leaf_194_clk channels.exp_counter\[1\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_127_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15916_ tt_um_rejunity_sn76489.chan\[0\].attenuation.in _07798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_155_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11039_ filters.sample_filtered\[1\] _03263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_95_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13691__A1 _05596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16896_ _00977_ _00843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_155_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15847_ _07598_ _07732_ _00646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_56_Left_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_91_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09647__B1 _01964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15778_ _07630_ _07682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17517_ _00587_ clknet_5_2__leaf_clk filters.high\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14729_ _06719_ _06722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11454__B1 _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17448_ _00518_ clknet_leaf_158_clk channels.accum\[3\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_172_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10009__A1 _02252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10096__I _01085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17379_ _00449_ clknet_leaf_131_clk channels.env_counter\[2\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_65_Left_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_93_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10980__A2 _03204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_151_Right_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_235_clk clknet_5_16__leaf_clk clknet_leaf_235_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_103_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11655__I _03039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09704_ channels.freq1\[12\] _02082_ _02077_ _02083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_74_Left_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09635_ channels.atk_dec3\[5\] _01991_ _01992_ channels.freq3\[13\] _02021_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_78_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09566_ channels.ch3_env\[2\] _01876_ _01886_ channels.freq1\[10\] _01955_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_136_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08517_ _01043_ _01008_ _01016_ _01044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_93_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11445__B1 _01420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09497_ channels.pw1\[0\] _01885_ _01887_ channels.freq1\[8\] _01888_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10799__A2 _03052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08861__A1 _01323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_83_Left_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10410_ _02669_ _02670_ _02671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_151_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11390_ _03566_ _01433_ _03572_ _00349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10341_ _02601_ _02602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13060_ _04918_ _05064_ _05065_ _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10272_ channels.env_vol\[0\]\[3\] channels.env_vol\[1\]\[3\] _02518_ _02533_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_143_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12011_ _04078_ _04079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_148_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_226_clk clknet_5_20__leaf_clk clknet_leaf_226_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_44_1195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11920__A1 _03534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_92_Left_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__15662__A2 _07592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16750_ _00867_ _00869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13962_ _05765_ _05845_ _05964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_161_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15701_ _07625_ _00607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12913_ _04470_ _04510_ _04919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16681_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[6\] _08399_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[6\]
+ _08424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13893_ _04642_ _05892_ _05895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16611__A1 _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15632_ _03391_ _07563_ _07564_ _03223_ _07565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_122_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12844_ _04703_ _04850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_122_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12779__A3 _04784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15563_ _03309_ _07488_ _07500_ _06066_ _07501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_12775_ _04780_ _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_17302_ _00372_ clknet_leaf_154_clk channels.accum\[1\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_173_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14514_ _06491_ _06492_ _06490_ _06510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11726_ channels.atk_dec3\[3\] _01439_ _03783_ channels.atk_dec2\[3\] _03817_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15494_ _07426_ _07432_ _07437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_16_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08852__A1 _01160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17233_ _00303_ clknet_leaf_172_clk channels.sample1\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14445_ _06440_ _06441_ _06442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11657_ _02687_ _03748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_126_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17164_ _00234_ clknet_leaf_144_clk channels.ctrl_reg3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10608_ _02562_ _02823_ _02867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14376_ _06236_ _06249_ _06374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11834__S1 _01170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11588_ _03689_ _03698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16115_ _07960_ _07892_ _07992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13327_ _05250_ _05333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_168_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17095_ _00165_ clknet_leaf_104_clk channels.ctrl_reg1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10539_ _02748_ _02749_ _02799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_51_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16046_ _07873_ _07919_ _07925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13258_ _05255_ _05263_ _05264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__17574__D _00644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_217_clk clknet_5_21__leaf_clk clknet_leaf_217_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_110_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12209_ _03239_ _03203_ _04189_ _04214_ _04215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__13900__A2 _05843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13189_ _05132_ _05192_ _05195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16948_ _00027_ clknet_leaf_239_clk channels.lfsr\[3\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11675__B1 _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14786__I _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16879_ _01189_ _00956_ _00965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16602__A1 _01319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09420_ _01812_ _01813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11770__S0 _01152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08784__I _01257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09351_ _01748_ _01749_ _01753_ _01754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_133_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09282_ _01706_ _01591_ _01710_ _01699_ _00099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08843__A1 _01300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_173_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14916__A1 filters.band\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13719__A2 _04403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10650__A1 _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10402__A1 _02662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10953__A2 _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14144__A2 _05690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_208_clk clknet_5_22__leaf_clk clknet_leaf_208_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_100_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10705__A2 _02777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09571__A2 _01954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08997_ _01449_ _01458_ _01459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11385__I _01089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13655__A1 _05568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_3_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09323__A2 _01734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09618_ channels.pw1\[4\] _02003_ _02004_ channels.ctrl_reg1\[4\] _02005_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_67_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10890_ _03126_ _03134_ _03140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_92_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_84_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11418__B1 _01568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09549_ channels.sus_rel2\[2\] _01936_ _01937_ channels.freq3\[2\] _01938_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_66_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12560_ _04226_ _04566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12630__A2 _04632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11511_ channels.pw1\[0\] _03643_ _03644_ _03645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12491_ _04410_ _04412_ _04497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_18_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14230_ _06216_ _06228_ _06229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_80_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14383__A2 _04632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15580__A1 channels.sample1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11442_ channels.accum\[1\]\[8\] _03602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_22_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14161_ _06103_ _06160_ _06161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11373_ channels.accum\[2\]\[3\] _03559_ _03562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10944__A2 _03080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10324_ _02577_ _02584_ _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13112_ _04535_ _04896_ _05118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__15476__B _07240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14092_ _04561_ _06086_ _06092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13043_ _04923_ _05049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10255_ _01306_ _02515_ _02516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_163_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_163_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10186_ _01533_ _02444_ _02445_ _02446_ _02447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__15990__I _02101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16802_ _00905_ _00907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_17782_ _00852_ clknet_leaf_200_clk channels.exp_periods\[0\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_156_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14994_ filters.filt_3 channels.sample3\[2\] _06965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16733_ _08463_ _08465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13945_ _05186_ _05947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_163_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11752__S0 _03832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16664_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[3\] _08398_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[3\]
+ _08410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13876_ _05772_ _05780_ _05878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_9_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15615_ _07538_ _07549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_147_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12827_ _04778_ _04786_ _04832_ _04833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_16595_ _08367_ _08369_ _08313_ _00757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_178_3680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_3691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15546_ filters.sample_buff\[3\] _07484_ _07485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12758_ _04211_ _04764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08825__A1 _01270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_155_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11709_ channels.atk_dec3\[5\] _01078_ _03780_ channels.atk_dec2\[5\] _01291_ channels.atk_dec1\[5\]
+ _03800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XTAP_TAPCELL_ROW_139_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_139_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15477_ _07419_ _07420_ _07421_ _07422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12689_ _04385_ _04695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_53_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17216_ _00286_ clknet_leaf_175_clk channels.sample2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_14428_ _06420_ _06424_ _06425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11807__S1 _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17147_ _00217_ clknet_leaf_144_clk channels.sus_rel2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_21_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14359_ _06356_ _04617_ _06357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15323__A1 _07277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17078_ _00148_ clknet_leaf_119_clk net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_123_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_139_Left_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16029_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\] _07909_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08920_ channels.freq3\[6\] _01076_ _01387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13885__A1 _05792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08851_ _01298_ _01323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_97_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_137_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_88_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08782_ _01102_ _01253_ _01256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_97_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_4__f_clk clknet_3_1_0_clk clknet_5_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_0_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15405__I _07355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_148_Left_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_177_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12860__A2 _04863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09403_ filters.mode_vol\[3\] _01794_ _01796_ _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_133_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10871__A1 _02029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09334_ channels.lfsr\[1\]\[22\] _01738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_62_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12612__A2 _04468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10623__A1 _02359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09265_ channels.lfsr\[3\]\[16\] _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_62_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_173_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09196_ _01635_ _01636_ _01628_ _01637_ _01605_ _01607_ _01638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__15562__A1 channels.sample3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_157_Left_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_71_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10926__A2 _01560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08689__I _01172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10040_ _02149_ _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_105_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11329__B _03517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11351__A2 _03534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13628__A1 _05630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12939__I _04858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11991_ _04043_ _04061_ _04062_ _00460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13730_ _05730_ _05733_ _05734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10942_ _03168_ _03052_ _03172_ _00301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12851__A2 _04855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13661_ _04562_ _05561_ _05574_ _05665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_42_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10873_ _03108_ _03121_ _03124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15400_ filters.low\[22\] _06836_ _07351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_27_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12612_ _04615_ _04468_ _04616_ _04617_ _04618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_16380_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[1\] _08192_ _08196_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13592_ _04220_ _04926_ _05597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_112_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15331_ _06919_ _07287_ _07288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_156_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12543_ _04356_ _04249_ _04357_ _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_66_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_156_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10090__A2 _02351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14356__A2 _04578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15262_ filters.high\[12\] _07062_ _07223_ _07224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15553__A1 channels.sample1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12474_ _04385_ _04480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_163_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_117_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17001_ _00080_ clknet_leaf_218_clk channels.lfsr\[2\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12367__A1 _04372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14213_ _05930_ _05075_ _06212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11425_ _03589_ _03591_ _01316_ _03592_ _00364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_15193_ _01771_ channels.sample3\[9\] _07157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_7 _01590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_134_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10917__A2 _03104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14144_ _04742_ _05690_ _06144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11356_ _03529_ _03531_ _03550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_162_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10393__A3 _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10307_ _01470_ _02541_ _02568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10922__I _02365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14075_ _05868_ _06075_ _05972_ _06076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11287_ _00999_ _01003_ _03493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13026_ _05028_ _05021_ _05032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10238_ _02484_ _02498_ _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_20_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10145__A3 channels.pw3\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09932__B _02243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10169_ _01284_ _02430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_179_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17765_ _00835_ clknet_leaf_82_clk tt_um_rejunity_sn76489.clk_counter\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09299__A1 _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14977_ _06939_ _05035_ _06948_ _06949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xrebuffer19 _05182_ net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_159_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16716_ _08449_ _08446_ _08452_ _00795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13928_ _05230_ _05930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_17696_ _00766_ clknet_leaf_223_clk channels.lfsr\[0\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16647_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[0\] _08263_ _08396_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10369__I _02543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10853__A1 channels.sample3\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13859_ _05856_ _05861_ _05862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_123_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16578_ _08314_ _08355_ _00754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15529_ _07462_ _07469_ _07470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09050_ channels.accum\[0\]\[15\] channels.accum\[1\]\[15\] channels.accum\[2\]\[15\]
+ channels.accum\[3\]\[15\] _00009_ _01153_ _01508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_44_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09952_ channels.freq3\[12\] _02258_ _02255_ _02259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_111_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08903_ _01337_ _01370_ _01371_ _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_09883_ _02209_ _02210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12530__A1 _04535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08834_ _01306_ _01307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16272__A2 _07742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12759__I _04764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08765_ channels.exp_counter\[2\]\[1\] _01090_ _01225_ _01241_ _01243_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_174_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_170_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08696_ channels.exp_periods\[2\]\[0\] _01180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_164_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14035__A1 _06030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09317_ _01650_ _01732_ _01733_ _01654_ _00111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_36_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09248_ channels.lfsr\[2\]\[15\] _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_111_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_201_clk_I clknet_5_23__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09179_ channels.lfsr\[1\]\[4\] _01623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_151_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_151_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11210_ filters.band\[12\] _03423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_160_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12190_ _04195_ _04196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_82_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput22 net22 bus_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_11141_ filters.sample_filtered\[8\] _03358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_216_clk_I clknet_5_21__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13849__A1 _05849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17048__CLK clknet_5_17__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11072_ filters.sample_filtered\[2\] _03276_ _03294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10023_ channels.atk_dec3\[7\] _02302_ _02303_ _02307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14900_ _06766_ _06877_ _06878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_15880_ _07754_ _07758_ _07761_ _07762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14831_ _06814_ _06815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_17550_ _00620_ clknet_leaf_5_clk filters.low\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14762_ _06735_ _06749_ _06750_ _06709_ _06751_ _06752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_11974_ channels.env_counter\[2\]\[8\] _04048_ _04049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_169_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_16501_ _08285_ _08290_ _08291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_158_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13713_ _05708_ _05716_ _05717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_58_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17481_ _00551_ clknet_leaf_32_clk filters.band\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10925_ _01321_ _03162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_158_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14693_ _06652_ _06685_ _06687_ _06688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__09978__I _02254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16432_ _08192_ _08233_ _08234_ _00729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09128__S1 _01304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13644_ _03251_ _03376_ _05648_ _05649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10856_ _03085_ _03103_ _03107_ _03108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16363_ _08176_ _08184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13575_ _05514_ _05580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_136_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10787_ _03037_ _03041_ _03042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_137_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15314_ _07271_ _07263_ _07264_ _07272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_171_3558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12526_ _04233_ _04245_ _04531_ _04532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__11260__A1 _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15526__A1 channels.sample1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16294_ _08144_ _00681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15245_ _07183_ _07207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_35_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12457_ _04383_ _04394_ _04463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_83_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11012__A1 _03204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11408_ channels.accum\[2\]\[17\] _01245_ _01530_ _01084_ _03583_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_15176_ _07095_ _07118_ _07140_ _07141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_12388_ _04387_ _04391_ _04393_ _04394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_50_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14127_ _06038_ _06039_ _06127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_11339_ _03532_ _03533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_123_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14058_ _05977_ _05979_ _06058_ _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__13304__A3 _05106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13009_ _05005_ _05013_ _05014_ _05015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_175_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11483__I _03624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14265__A1 _04644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08550_ clk_ctr\[0\] _01066_ _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17748_ _00818_ clknet_leaf_55_clk tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__16495__B _08244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08481_ _01002_ _01003_ _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14017__A1 _06015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17679_ _00749_ clknet_leaf_68_clk tt_um_rejunity_sn76489.tone\[1\].gen.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08495__A2 _01022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12579__A1 _04583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09444__A1 channels.ctrl_reg2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09102_ _01536_ _01543_ _01553_ _01554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_174_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08798__A3 _01082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_143_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14743__B _06734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09033_ channels.freq3\[14\] _01080_ _01492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_96_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14740__A2 _06731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_74_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09935_ _02208_ _01833_ _02246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_0_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09866_ _02188_ _02194_ _02198_ _00199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_70_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08817_ _01289_ _01290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09797_ _02131_ _02142_ _02148_ _00180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13059__A2 _04221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_82_clk_I clknet_5_9__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08748_ _01229_ _00046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_36_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09683__A1 filters.cutoff_lut\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14008__A1 _04487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08679_ _01162_ _01163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_95_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09683__B2 channels.ch3_env\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09798__I _01017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10710_ _02960_ _02966_ _02967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11490__A1 channels.freq1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15756__A1 _03411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11690_ channels.sus_rel3\[0\] _01439_ _03780_ channels.sus_rel2\[0\] _03781_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_67_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_97_clk_I clknet_5_13__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10641_ _02897_ _02898_ _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_36_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13231__A2 _04371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_153_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16852__C _01069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13360_ _05258_ _05261_ _05366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_1_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10572_ channels.sample3\[1\] _02784_ _02832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_165_Right_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__17667__D _00737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_20_clk_I clknet_5_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12311_ _04316_ _04317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_114_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09747__B _02113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13291_ _05265_ _05297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_51_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15030_ _06969_ _06998_ _06999_ _07000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_107_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12242_ _04233_ _04245_ _04248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_133_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_155_clk_I clknet_5_29__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12173_ _04178_ _04179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_82_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11124_ filters.sample_filtered\[7\] _03342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_16981_ _00060_ clknet_leaf_180_clk channels.accum\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13783__I _05700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13298__A2 _05216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14495__A1 _06305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15932_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[1\] _07809_ _07814_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_11055_ _03267_ _03261_ _03277_ _03278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10006_ channels.atk_dec3\[1\] _02292_ _02294_ _02296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15863_ tt_um_rejunity_sn76489.chan\[2\].attenuation.in _07745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_129_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14247__A1 _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17602_ _00672_ clknet_leaf_41_clk spi_dac_i.spi_dat_buff_0\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14814_ _06753_ _06797_ _06799_ _06800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_157_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15794_ _07630_ _07694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_118_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17533_ _00603_ clknet_leaf_82_clk filters.sample_buff\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_14745_ _06732_ _06736_ _06737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_171_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11957_ channels.env_counter\[2\]\[5\] _04030_ _04035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09674__A1 channels.atk_dec1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10284__A2 _02543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17464_ _00534_ clknet_leaf_2_clk filters.band\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10908_ channels.sample2\[5\] _03150_ _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14676_ _06583_ _06587_ _06671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15747__A1 _07659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_103_Left_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11888_ _03947_ _03968_ _03973_ _03974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_16415_ _08219_ _08221_ _08222_ _00724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_27_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13627_ _03332_ _04522_ _05487_ _05632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_17395_ _00465_ clknet_leaf_132_clk channels.env_counter\[1\]\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_108_clk_I clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10839_ _03064_ _03069_ _03067_ _03092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16346_ _08173_ _00704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13558_ _04562_ _05563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_109_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_132_Right_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11784__A2 _03874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12509_ _04503_ _04514_ _04515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_16277_ _08135_ _08136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13489_ _05341_ _05495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_89_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15228_ _07190_ _05646_ _07191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_140_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14722__A2 _06714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15159_ _07105_ _07110_ _07124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_1_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_112_Left_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14789__I _06689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09720_ _02093_ _02094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_52_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09651_ _01934_ net27 _02036_ _02037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14238__A1 filters.band\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08602_ channels.lfsr\[3\]\[5\] _01112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09582_ _01886_ _01970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_136_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08533_ _01040_ _01030_ _01025_ _01056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_54_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09665__A1 channels.freq1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09665__B2 channels.pw3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13461__A2 _04182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15738__A1 _03329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09411__I _01006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09417__A1 _01807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09968__A2 _02266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09016_ _01468_ _01470_ _01476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14713__A2 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12724__A1 _04728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11388__I _02974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12724__B2 _04259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14477__A1 _06472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09918_ _02215_ _02227_ _02233_ _00216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_146_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09849_ _02185_ _02181_ _02186_ _00194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_154_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12860_ _04859_ _04863_ _04865_ _04866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_107_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11811_ _03803_ _03857_ _03826_ _03884_ _03902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_69_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12791_ _04792_ _04796_ _04797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_96_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14530_ _06524_ _06525_ _06526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11742_ channels.env_counter\[0\]\[2\] channels.env_counter\[1\]\[2\] channels.env_counter\[2\]\[2\]
+ channels.env_counter\[3\]\[2\] _03832_ _01171_ _03833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_95_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09321__I _01730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14461_ _06454_ _06455_ _06457_ _06458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_166_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11673_ _02711_ _03539_ _03763_ _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14401__A1 _03361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16200_ _07834_ _08073_ _08074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_12_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13412_ _04874_ _04951_ _05418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_14_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17180_ _00250_ clknet_leaf_76_clk channels.sus_rel3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10624_ _02358_ _02882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14392_ _06305_ _06389_ _06390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14952__A2 channels.sample3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16131_ _07977_ _08005_ _08006_ _08007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13343_ _04198_ _04926_ _05349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10555_ _02809_ _02814_ _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_180_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16062_ _07823_ _07827_ _07817_ _07910_ _07941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_13274_ _05279_ _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13507__A3 _04758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10486_ _02629_ _02745_ _02746_ _02747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_122_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15013_ _06982_ _06983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_12225_ _04230_ _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_20_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12156_ _03190_ _03312_ _03196_ filters.high\[5\] _04162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_TAPCELL_ROW_166_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_166_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11107_ filters.sample_filtered\[6\] _03326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_12087_ _04061_ _04119_ _04124_ _00494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16964_ _00043_ clknet_leaf_211_clk channels.env_vol\[3\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15915_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[1\] _07797_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_11038_ _03213_ _03260_ _03262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09895__A1 _02215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16895_ _00962_ channels.exp_periods\[1\]\[1\] _00975_ _00977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13691__A2 _05597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15846_ spi_dac_i.counter\[1\] _07728_ _07731_ _07732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09647__A1 filters.bp vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12989_ _04503_ _04514_ _04995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_15777_ _06783_ _07677_ _07681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09647__B2 channels.sus_rel1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17516_ _00586_ clknet_5_1__leaf_clk filters.high\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14728_ _06720_ _06712_ _06721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14659_ _06542_ _06558_ _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_17447_ _00517_ clknet_leaf_162_clk channels.accum\[3\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_180_clk clknet_5_19__leaf_clk clknet_leaf_180_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_27_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17378_ _00448_ clknet_leaf_204_clk channels.env_vol\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_160_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_31_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16329_ channels.env_vol\[1\]\[3\] _08160_ _08164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_120_Left_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09583__B1 _01970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09406__I _01800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09703_ _02073_ _02082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_96_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09886__A1 _02179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09634_ channels.sus_rel3\[5\] _01963_ _01970_ channels.freq1\[13\] _02020_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_179_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09565_ _01855_ _01954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09638__A1 channels.pw2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09638__B2 channels.freq2\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08516_ _01042_ _01043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_172_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09496_ _01886_ _01887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_33_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_102_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_171_clk clknet_5_24__leaf_clk clknet_leaf_171_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_163_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13198__A1 _05142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09810__A1 channels.sus_rel1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10340_ _02583_ _02601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14698__A1 _06599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14931__B _06775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12007__I _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10271_ _01143_ channels.env_vol\[3\]\[3\] _02531_ _02532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_12010_ _04077_ _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_148_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11846__I _03936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11920__A2 _04002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13961_ _05879_ _05962_ _05963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__11067__B _03288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12912_ _04229_ _04483_ _04918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_15700_ channels.exp_periods\[3\]\[2\] _07625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16680_ _08419_ _08423_ _00788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10487__A2 _02543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13892_ _05795_ _05797_ _05893_ _05894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_159_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12843_ _04847_ _04269_ _04181_ _04848_ _04849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_15631_ _02029_ _07549_ _07564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09629__A1 _02008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12228__A3 _04221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_122_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15562_ channels.sample3\[4\] _07453_ _07500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12774_ _04779_ _04780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_68_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09051__I _01508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14513_ _06491_ _06492_ _06490_ _06509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_83_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17301_ _00371_ clknet_leaf_169_clk channels.accum\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11725_ _03803_ _03815_ _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_15493_ filters.high\[31\] _07436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_56_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_162_clk clknet_5_25__leaf_clk clknet_leaf_162_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_127_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14444_ _04318_ _05585_ _06441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17232_ _00302_ clknet_leaf_172_clk channels.sample1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08890__I _01257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11656_ _02721_ _03747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_83_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12936__A1 _04863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17163_ _00233_ clknet_leaf_144_clk channels.ctrl_reg3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10607_ _02810_ _02813_ _02865_ _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14375_ _06263_ _06264_ _06267_ _06373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__10925__I _01321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11587_ _03695_ _03697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16114_ _07800_ _07990_ _07991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_135_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13326_ _05331_ _05321_ _05332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_107_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17094_ _00164_ clknet_leaf_110_clk channels.ctrl_reg1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10538_ _02748_ _02749_ _02798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_168_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16045_ _07869_ _07924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13257_ _05257_ _05262_ _05263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__16612__I _08374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10469_ _02693_ _02727_ _02729_ _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_122_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12208_ filters.high\[0\] _04214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_13188_ _05058_ _05086_ _05095_ _05194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_12139_ _04151_ _00519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16947_ _00026_ clknet_leaf_238_clk channels.lfsr\[3\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09868__A1 channels.ctrl_reg2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14861__A1 _06761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11675__A1 channels.sus_rel2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11675__B2 channels.sus_rel1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16878_ _00940_ _00954_ _00964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__11770__S1 _01171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15829_ _07598_ _07716_ _00644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_176_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14613__A1 _06403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09350_ _01752_ _01753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_75_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_47_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09281_ _01707_ _01708_ _01701_ _01709_ _01679_ _01680_ _01710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_30_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16366__A1 _03964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15169__A2 _07133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_153_clk clknet_5_29__leaf_clk clknet_leaf_153_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_7_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09896__I _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10650__A2 _02823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14916__A2 _03476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13719__A3 _04805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_5_19__f_clk_I clknet_3_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08996_ _01456_ _01457_ _01458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_103_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09136__I _01584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_143_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_3_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09617_ _01941_ _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_67_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09548_ _01870_ _01937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_84_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_148_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09479_ _01832_ _01860_ _01870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_144_clk clknet_5_30__leaf_clk clknet_leaf_144_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__16357__A1 channels.ch3_env\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11510_ _03516_ _03644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_114_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12490_ _04462_ _04465_ _04495_ _04496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_47_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11441_ _03600_ _01406_ _03601_ _00371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_22_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14160_ _06136_ _06159_ _06160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11372_ _03561_ _03557_ _01348_ _03558_ _00342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_150_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13111_ _04901_ _04904_ _05116_ _05117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_46_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10323_ _02524_ _02543_ _02583_ _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_14091_ _06004_ _06020_ _06090_ _06091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15332__A2 _07033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13343__A1 _04198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13042_ _05044_ _05047_ _05048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_10254_ channels.ch3_env\[2\] _02515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11354__B1 _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_163_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_163_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10185_ channels.pw1\[6\] _02430_ _02446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_180_3730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16801_ _00905_ _00906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17781_ _00851_ clknet_leaf_206_clk channels.exp_counter\[3\]\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14993_ _06962_ _06963_ _06964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__14843__A1 _06720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16732_ _08463_ _08464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13944_ _05941_ _05945_ _05946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__11752__S1 _03842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16596__A1 _08242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16663_ _08408_ _08409_ _00785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13875_ _05432_ _05871_ _05872_ _05876_ _05877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_15614_ filters.sample_buff\[7\] _07543_ _07548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12200__I _04182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12826_ _04782_ _04785_ _04832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_57_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16594_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[8\] _08274_ _08368_ _08369_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_69_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_178_3681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_3692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15545_ _07446_ _07484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12757_ _04287_ _04505_ _04763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_135_clk clknet_5_31__leaf_clk clknet_leaf_135_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_29_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11708_ _03788_ _03798_ _03532_ _03799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_15476_ _07419_ _07420_ _07240_ _07421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_139_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12688_ _04467_ _04694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_112_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12909__A1 _04855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14427_ _06421_ _06422_ _06423_ _06424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_4_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17215_ _00285_ clknet_leaf_179_clk channels.sample2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_86_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11639_ _01750_ _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_25_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12385__A2 _04390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17146_ _00216_ clknet_leaf_123_clk channels.sus_rel2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_141_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14358_ filters.band\[28\] _06356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13309_ _04267_ _04179_ _04781_ _04803_ _05315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_17077_ _00147_ clknet_leaf_125_clk net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__16520__A1 _08274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14289_ _06287_ _06179_ _06288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_97_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13334__A1 _04254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09538__B1 _01905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16028_ _07819_ _07907_ _07908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_110_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08850_ _01321_ _01322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_88_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08781_ _01254_ _01255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_88_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14797__I _06760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09402_ _01767_ _01793_ _01798_ _00135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_88_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09333_ _01715_ _01722_ _01726_ _01718_ _00123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_158_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12612__A3 _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09264_ channels.lfsr\[1\]\[16\] _01696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10623__A2 _02880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15011__A1 _04158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09195_ channels.lfsr\[3\]\[6\] _01637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10139__A1 channels.pw1\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11351__A3 _03544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08979_ _01440_ _01441_ _01442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__13628__A2 _05631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11990_ channels.env_counter\[2\]\[11\] _04048_ _04062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10941_ channels.sample1\[6\] _03170_ _03172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16578__A1 _08314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12851__A3 _04856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12020__I _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13660_ _04645_ _05663_ _05572_ _05664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_39_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10862__A2 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10872_ _03054_ _03122_ _03123_ _00280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12611_ _04599_ _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_117_clk clknet_5_27__leaf_clk clknet_leaf_117_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_27_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13591_ _04236_ _04861_ _05596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_109_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15330_ _07284_ _07286_ _07287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_12542_ _04533_ _04534_ _04547_ _04548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_156_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15261_ _03721_ _07223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12473_ _04236_ _04278_ _04479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14212_ _05465_ _05049_ _06211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_17000_ _00079_ clknet_leaf_212_clk channels.lfsr\[2\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13564__A1 _04630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11424_ _01101_ _03592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15192_ _07153_ _07154_ _07155_ _07156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09232__A2 _01659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_8 _01590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14143_ _04529_ _06008_ _06143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11355_ _03547_ _03548_ _03549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_85_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10306_ _02539_ _02567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_14074_ _05856_ _05861_ _06075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11286_ net12 _03492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13025_ _05017_ _05030_ _05031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_123_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10237_ _02486_ _02494_ _02497_ _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_10168_ _02426_ _02428_ channels.pw3\[7\] _02429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__10550__A1 _02522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17764_ _00834_ clknet_leaf_81_clk tt_um_rejunity_sn76489.clk_counter\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09299__A2 _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14976_ filters.low\[2\] _06947_ _06948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10099_ _02359_ _02361_ _02362_ _00268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16715_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[5\] _08447_ _08451_ _08452_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13927_ _04752_ _05229_ _05929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17695_ _00765_ clknet_leaf_219_clk channels.lfsr\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10302__A1 _02555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_179_Right_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16646_ _08267_ _08394_ _08395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13858_ _05857_ _05859_ _05860_ _05861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_69_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12809_ _04787_ _04798_ _04815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_44_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16577_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[5\] _08347_ _08353_ _08354_
+ _08355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xclkbuf_leaf_108_clk clknet_5_15__leaf_clk clknet_leaf_108_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_130_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13789_ _05708_ _05716_ _05791_ _05792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_32_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15528_ filters.sample_buff\[1\] _07468_ _07469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_57_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15459_ _07388_ _07404_ _07405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_170_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17129_ _00199_ clknet_leaf_118_clk channels.ctrl_reg2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_52_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09951_ _02246_ _02258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_110_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08902_ _01364_ _01369_ _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_148_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09882_ _02208_ _01838_ _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_110_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08734__A1 _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08833_ _01305_ _01306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12530__A2 _04171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08764_ _01242_ _00049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09414__I _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11165__B _03380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08695_ _01178_ _01179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_146_Right_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10844__A2 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12775__I _04780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09316_ _01645_ _01732_ _01733_ _01648_ _00110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_76_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13794__A1 _04487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12597__A2 _04297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09247_ _01675_ _01659_ _01681_ _01674_ _00093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10295__I channels.ch3_env\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09178_ channels.lfsr\[0\]\[4\] _01622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_90_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_79_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_151_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_151_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput23 net23 bus_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_11140_ _03342_ _03327_ _03328_ _03357_ _00314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_31_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_112_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11071_ _03292_ _03293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_101_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10022_ _02240_ _02301_ _02306_ _00247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14830_ _06777_ _06813_ _06814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_11973_ _04011_ _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14761_ _06731_ _06741_ _06734_ _06751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_86_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16500_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[4\] _08269_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[4\]
+ _08290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_58_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13712_ _05711_ _05715_ _05716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10924_ _03160_ _03141_ _03161_ _00294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_158_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14692_ _06512_ _06598_ _06686_ _06687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17480_ _00550_ clknet_leaf_23_clk filters.band\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_158_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_113_Right_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16431_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[14\] _08192_ _08195_ _08234_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_116_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10855_ _03086_ _03102_ _03107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13643_ _05647_ _03219_ _05648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_175_3640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13574_ _05494_ _05524_ _05578_ _05579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_54_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16362_ _03958_ _08177_ _08183_ _00710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_137_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10786_ _03038_ _03040_ _03041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_9_clk_I clknet_5_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_136_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12525_ _04530_ _04193_ _04202_ _04531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_15313_ _07246_ _07249_ _07271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_TAPCELL_ROW_171_3559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16293_ channels.env_counter\[3\]\[2\] _08144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_136_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11260__A2 _03194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16723__A1 _08456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17762__CLK clknet_5_9__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12456_ _04448_ _04461_ _04462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_15244_ _07179_ _07204_ _07205_ _07206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_23_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_10_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11407_ _03580_ _03581_ _01524_ _03582_ _00356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_112_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15175_ _07113_ _07117_ _07140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11012__A2 _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12387_ _04392_ _04280_ _04393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14126_ _06038_ _06039_ _06126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11338_ _03530_ _03531_ _03532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_22_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14057_ _05997_ _06000_ _06057_ _06058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_11269_ _03467_ _03236_ _03469_ _03478_ _03479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__16620__I _08380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_176_Left_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13008_ _05011_ _05012_ _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_94_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11720__C2 channels.atk_dec1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14265__A2 _06261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17747_ _00817_ clknet_5_8__leaf_clk tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12276__A1 _04281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14959_ _06909_ _06931_ _06932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09141__A1 _01043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08480_ net17 _01010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_17678_ _00748_ clknet_leaf_56_clk tt_um_rejunity_sn76489.chan\[2\].attenuation.in
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14017__A2 _06016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_7_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16629_ _01673_ _08386_ _08387_ _01676_ _00773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_169_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09444__A2 _01830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09101_ _01549_ _01553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_143_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15517__A2 _07458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09032_ _01490_ _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08955__A1 _01337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09934_ _02104_ _02245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_74_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09865_ channels.ctrl_reg2\[2\] _02195_ _02189_ _02198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_175_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08816_ _01288_ _01289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09796_ channels.sus_rel1\[3\] _02143_ _02146_ _02148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13059__A3 _04274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17635__CLK clknet_5_23__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08747_ channels.exp_counter\[1\]\[2\] _01105_ _01228_ _01220_ _01229_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08678_ _01161_ _01162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_96_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14008__A2 _06008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13767__A1 _05686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10640_ _02851_ _02854_ _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10571_ _02788_ _02830_ _02831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_10_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12310_ _04315_ _04316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_23_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13290_ _05203_ _05241_ _05296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_107_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12241_ _04183_ _04193_ _04202_ _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_106_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_131_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12172_ _03331_ _04177_ _04178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_20_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11123_ _03326_ _03327_ _03328_ _03341_ _00313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_16980_ _00059_ clknet_leaf_186_clk channels.accum\[0\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_102_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15931_ _07812_ _07813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11054_ filters.sample_filtered\[2\] _03276_ _03277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10505__A1 _02662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10005_ _02245_ _02291_ _02295_ _00241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_15862_ _04170_ _07743_ _07744_ _07710_ _00649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_129_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14247__A2 _05891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17601_ _00671_ clknet_leaf_41_clk spi_dac_i.spi_dat_buff_0\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14813_ _06779_ _06780_ _06788_ _06798_ _06799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_15793_ _06818_ _07690_ _07693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09123__A1 _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09989__I _02254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17532_ _00602_ clknet_leaf_82_clk filters.sample_buff\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_114_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14744_ net30 _06733_ _06735_ _06736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11956_ _04009_ _04032_ _04033_ _04034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_58_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17463_ _00533_ clknet_leaf_1_clk filters.band\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15005__B _06952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10928__I _01460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10907_ _03147_ _02973_ _03151_ _00287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_169_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14675_ _05268_ _05626_ _06670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10284__A3 _02544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11887_ _03970_ _03972_ _03947_ _03973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_157_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16414_ _08194_ _08222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_129_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13626_ _03316_ _04163_ _05208_ _05631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_10838_ _03087_ _03089_ _03090_ _03091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_17394_ _00464_ clknet_leaf_132_clk channels.env_counter\[1\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_15_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16345_ _01228_ _01317_ _01258_ channels.exp_counter\[0\]\[2\] _08173_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09938__B _02243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13557_ _05560_ _05561_ _05451_ _05562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__16615__I _08382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10769_ _02999_ _03004_ _03024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12508_ _04509_ _04513_ _04514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_54_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16276_ _03940_ _08135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13488_ _05461_ _05493_ _05494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_180_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12439_ _04444_ _04445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15227_ _07188_ _07189_ _07190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_39_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15158_ _07105_ _07110_ _07123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10744__A1 _02710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13974__I _05543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14109_ _06033_ _06034_ _06108_ _06109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_91_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15089_ _03310_ _07022_ _07057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11708__B _03532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11494__I _03624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09362__A1 _01762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09650_ _01808_ _02036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14238__A2 _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08601_ _01111_ _00017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_145_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_200_clk_I clknet_5_23__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09581_ channels.ch3_env\[3\] _01877_ _01885_ channels.pw1\[3\] _01969_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_145_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08532_ _01016_ _00130_ _01055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13997__A1 _05905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13214__I _04780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_215_clk_I clknet_5_21__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_98_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_30_clk clknet_5_0__leaf_clk clknet_leaf_30_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_45_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09015_ _01463_ _01409_ _01475_ _01421_ _00067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_76_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08928__A1 _01337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16260__I _07741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09917_ channels.sus_rel2\[3\] _02228_ _02232_ _02233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12488__A1 _04475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_97_clk clknet_5_13__leaf_clk clknet_leaf_97_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09848_ channels.pw2\[9\] _02182_ _02176_ _02186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_146_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09779_ _01807_ _02133_ _02136_ _00174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_73_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11810_ _03857_ _03897_ _03900_ _03901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_68_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12790_ _04793_ _04794_ _04795_ _04796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_0_139_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09656__A2 _02038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output28_I net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11741_ _03831_ _03832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_68_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11672_ channels.sus_rel3\[4\] _01081_ _01281_ channels.sus_rel2\[4\] _03762_ _03763_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_7_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14460_ _06456_ _04617_ _06457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_165_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14401__A2 _06397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13411_ _05413_ _05409_ _05417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_48_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10623_ _02359_ _02880_ _02881_ _00273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_12_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14391_ _06308_ _06388_ _06389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09758__B _02120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_21_clk clknet_5_3__leaf_clk clknet_leaf_21_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_107_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16130_ _07981_ _08002_ _08006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_24_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13342_ _04265_ _05347_ _05348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10554_ _02810_ _02813_ _02814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_10_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16061_ _07910_ _07940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13273_ _05077_ _05279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_121_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10485_ _02631_ _02639_ _02746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__13507__A4 _04946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13912__A1 _04451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12224_ _04229_ _04230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15012_ _06981_ _06982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_121_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09592__A1 channels.ctrl_reg2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09592__B2 channels.ctrl_reg3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12155_ _04160_ _04161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_166_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_166_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11106_ _03309_ _03265_ _03266_ _03325_ _00312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_12086_ channels.env_counter\[0\]\[11\] _04120_ _04124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16963_ _00042_ clknet_leaf_211_clk channels.env_vol\[3\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_88_clk clknet_5_12__leaf_clk clknet_leaf_88_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15914_ _07792_ _07794_ _07795_ _07796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_21_1164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13140__A2 _05145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11037_ _03213_ _03260_ _03261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_16894_ _00976_ _00842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15845_ spi_dac_i.counter\[1\] _07729_ _07730_ _07731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_8_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15776_ _06774_ _07640_ _07680_ _00627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12988_ _04512_ _04642_ _04509_ _04994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_59_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17515_ _00585_ clknet_leaf_37_clk filters.high\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14727_ _06719_ _06720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11939_ _03833_ _04015_ _04020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_115_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_157_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_129_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17446_ _00516_ clknet_leaf_151_clk channels.accum\[3\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08950__S0 _01148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14658_ _06614_ _05982_ _06653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13609_ _05611_ _05612_ _05613_ _05614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_7_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17377_ _00447_ clknet_leaf_214_clk channels.env_vol\[0\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14589_ _04924_ _05626_ _06585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_31_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16328_ _03954_ _08158_ _08163_ _00696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_171_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_153_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_81_clk_I clknet_5_9__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16259_ _08121_ _08124_ _00666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_129_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09583__A1 channels.pw3\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09583__B2 channels.freq1\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11390__A1 _03566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15656__A1 filters.sample_buff\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_96_clk_I clknet_5_13__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_79_clk clknet_5_12__leaf_clk clknet_leaf_79_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09702_ _02073_ _02081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09633_ filters.cutoff_lut\[14\] _01988_ _02019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_179_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09564_ channels.pw3\[10\] _01842_ _01848_ channels.pw2\[2\] _01952_ _01953_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_136_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_69_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_1__f_clk_I clknet_3_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08515_ net17 _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_clkbuf_leaf_154_clk_I clknet_5_29__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09495_ _01854_ _01846_ _01886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12642__A1 filters.res_lut\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_34_clk_I clknet_5_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_65_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13198__A2 _05147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_169_clk_I clknet_5_24__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_49_clk_I clknet_5_10__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14698__A2 _06601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10270_ _01305_ _02530_ _02531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_108_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09574__A1 _01933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_107_clk_I clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13960_ _05882_ _05961_ _05962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__11067__C _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11133__A1 _03345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12911_ _04853_ _04915_ _04916_ _04917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_161_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13891_ _04597_ _05892_ _05798_ _05893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10487__A3 _02638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12881__A1 _03302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11684__A2 _03535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11862__I _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15630_ _07549_ _07563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12842_ _04237_ _04848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_158_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16874__B _00940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15561_ filters.sample_buff\[3\] _07493_ _07499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12773_ filters.cutoff_lut\[13\] _04442_ _04779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_84_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17300_ _00370_ clknet_leaf_188_clk channels.accum\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14512_ _05544_ _06508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_167_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11724_ _03805_ _03814_ _03815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_139_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15492_ _07424_ _07434_ _07435_ _00588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_166_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14386__A1 _05563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17231_ _00301_ clknet_leaf_170_clk channels.sample1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_182_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12693__I _04255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14443_ _04453_ _05500_ _06440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11655_ _03039_ _03746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_153_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17162_ _00232_ clknet_5_26__leaf_clk channels.pw3\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_24_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10606_ _02811_ _02812_ _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_11586_ _03695_ _03696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14374_ _06311_ _06371_ _06372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_181_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16113_ _07882_ _07989_ _07990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_13325_ _05323_ _05330_ _05331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10537_ _02795_ _02761_ _02796_ _02797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17093_ _00163_ clknet_leaf_110_clk channels.ctrl_reg1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_168_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15886__A1 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[2\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14689__A2 _06682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16044_ _07597_ _07923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13256_ _05258_ _05261_ _05262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10468_ _02683_ _02693_ _02694_ _02728_ _02729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_150_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12207_ _04172_ _04210_ _04212_ _04213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_161_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13187_ _05132_ _05192_ _05193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10399_ _02656_ _02658_ _02660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_86_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11372__B2 _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12138_ channels.accum\[3\]\[17\] _04151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12069_ _04106_ _04114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_159_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16946_ _00025_ clknet_leaf_236_clk channels.lfsr\[3\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_8_Left_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_1_clk clknet_5_4__leaf_clk clknet_leaf_1_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_159_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12872__A1 _04821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16877_ _01208_ _00938_ _00963_ _00838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_95_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15828_ _07443_ _07714_ _07716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_35_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11427__A2 _03593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15759_ _06714_ _07632_ _07668_ _00622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09280_ channels.lfsr\[3\]\[19\] _01709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08923__S0 _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17429_ _00499_ clknet_leaf_164_clk channels.adsr_state\[2\]\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14129__A1 _04376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11168__B _03383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08995_ _01450_ _01447_ _01455_ _01457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_103_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13104__A2 _04163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14301__A1 _06168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11115__A1 _03329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12778__I _04783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09616_ _01884_ _02003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_104_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14604__A2 _03377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09547_ _01868_ _01936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_84_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09478_ _01868_ _01869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_4_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11631__B _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11440_ channels.accum\[1\]\[7\] _03593_ _03601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10929__A1 channels.sample1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09795__A1 _02112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11371_ channels.accum\[2\]\[2\] _03561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13110_ _04902_ _04903_ _05116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_33_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10322_ _01688_ _02580_ _02582_ _02583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_14090_ _06002_ _06021_ _06090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_81_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11729__I0 channels.atk_dec1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13041_ _04952_ _04991_ _05014_ _05046_ _04993_ _05047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_10253_ _02513_ _02514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13343__A2 _04926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_29__f_clk clknet_3_7_0_clk clknet_5_29__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11354__A1 channels.ctrl_reg3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09327__I _01730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11354__B2 channels.ctrl_reg1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10184_ _02426_ _02405_ channels.pw3\[6\] _02445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__15773__B _07671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_180_3720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16800_ _00879_ _00904_ _00905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__15096__A2 _07061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_180_3731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08770__A2 _01245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17780_ _00850_ clknet_leaf_197_clk channels.exp_counter\[3\]\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14992_ filters.filt_1 channels.sample1\[2\] channels.sample2\[2\] filters.filt_2
+ _06963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12449__A4 _04453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16731_ _08461_ _08462_ _08444_ _08463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_13943_ _05942_ _05944_ _05945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_88_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16662_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[2\] _08345_ _08339_ _08409_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13874_ _05873_ _05874_ _05875_ _05876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_69_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15613_ _07536_ _07547_ _07435_ _00597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_12825_ _04793_ _04829_ _04830_ _04831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_16593_ _08238_ _08362_ _08366_ _08368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_178_3682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10001__I _02290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_178_3693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15544_ _07382_ _07483_ _00592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_96_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12756_ _04749_ _04761_ _04762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10093__A1 _01070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11707_ channels.atk_dec1\[1\] channels.sus_rel1\[1\] _03784_ _03798_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_166_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15475_ _07408_ _07412_ _07411_ _07420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_56_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12687_ _04520_ _04692_ _04693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_72_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15020__A2 channels.sample3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17214_ _00284_ clknet_leaf_179_clk channels.sample2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_154_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14426_ _04819_ _05075_ _06423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12909__A2 _04856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11638_ _03731_ _03732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_170_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_170_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17145_ _00215_ clknet_leaf_124_clk channels.sus_rel2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14357_ _04600_ _06093_ _06355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11569_ channels.freq3\[2\] _03681_ _03682_ _03685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11593__A1 channels.pw3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13308_ _04273_ _04800_ _05314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17076_ _00146_ clknet_leaf_119_clk net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14288_ _06176_ _06287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09538__A1 _01927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16027_ _07904_ _07906_ _07907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09538__B2 clk_trg\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13239_ _05157_ _05163_ _05245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_62_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08780_ _01253_ _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_127_Right_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13098__A1 _03270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16929_ _08449_ _00993_ _00995_ _00858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_137_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12845__A1 _04848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09710__A1 _01814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09401_ filters.mode_vol\[2\] _01794_ _01796_ _01798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_87_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09332_ _01710_ _01722_ _01726_ _01713_ _00122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_62_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13270__A1 _05184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12612__A4 _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09263_ channels.lfsr\[0\]\[16\] _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15011__A2 _04776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09194_ channels.lfsr\[1\]\[6\] _01636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_132_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09777__A1 _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11584__A1 _03677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15078__A2 channels.sample1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08978_ channels.freq2\[10\] _01278_ _01290_ channels.freq1\[10\] _01441_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__13628__A3 _05632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09701__A1 _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10940_ _03168_ _03013_ _03171_ _00300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14589__A1 _04924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16708__I _08445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10871_ _02029_ _03105_ _03123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15250__A2 channels.sample2\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12610_ _04578_ _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_27_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13590_ _04476_ _05077_ _05595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_151_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10075__A1 _02324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12541_ _04545_ _04546_ _04547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_26_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_156_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15260_ _07203_ _07221_ _07222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_152_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12472_ _04477_ _04476_ _04478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_173_3590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14211_ _06204_ _06209_ _06210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_108_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11423_ _03590_ _03591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14761__A1 _06731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09766__B _02120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15191_ _07130_ _07131_ _07155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_34_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10378__A2 _02569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_9 _01590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_134_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11354_ channels.ctrl_reg3\[0\] _01581_ _01295_ channels.ctrl_reg1\[0\] _03548_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_132_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14142_ _06048_ _06140_ _06141_ _06142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_61_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_89_Left_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10305_ _02506_ _02564_ _02565_ _02566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_11285_ net13 _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_14073_ _03299_ _06073_ _05968_ _05970_ _06074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_123_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10236_ _01266_ channels.ctrl_reg3\[6\] channels.ctrl_reg1\[6\] _01252_ _02496_ _02497_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_13024_ _05021_ _05028_ _05029_ _05030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_158_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08743__A2 _01105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10167_ _02427_ _02428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10550__A2 _02622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17763_ _00833_ clknet_leaf_86_clk tt_um_rejunity_sn76489.clk_counter\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14975_ _06944_ _06946_ _06947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10098_ channels.sync_outs\[2\] _01245_ _02362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16714_ _08450_ _08451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13926_ _04801_ _05183_ _05928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17694_ _00764_ clknet_leaf_220_clk channels.lfsr\[0\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_98_Left_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16645_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[0\] _08393_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[0\]
+ _08394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_16_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13857_ _05752_ _05755_ _05860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12808_ _04811_ net50 _04813_ _04814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_44_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16576_ _08349_ _08352_ _08301_ _08354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13252__A1 _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13788_ _05710_ _05790_ _05715_ _05791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_44_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10066__A1 _02316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_174_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15527_ _07466_ _07467_ _07468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_12739_ _04732_ _04736_ _04744_ _04745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_72_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_155_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15458_ _07386_ _07398_ _07404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_182_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11698__S _03784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09759__A1 _01819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14409_ _06404_ _06405_ _06406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14752__A1 _06722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15389_ _07321_ _07336_ _07340_ _07341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11566__A1 _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17128_ _00198_ clknet_5_27__leaf_clk channels.ctrl_reg2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_13_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14504__A1 _03380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09950_ _02246_ _02257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17059_ _00129_ clknet_leaf_94_clk filters.res_filt\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_3_3_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08901_ _01364_ _01369_ _01370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09881_ _01779_ _02208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_5_12__f_clk clknet_3_3_0_clk clknet_5_12__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_57_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08832_ _01142_ _01305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_100_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08763_ channels.exp_counter\[2\]\[0\] _01090_ _01218_ _01241_ _01242_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_139_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15480__A2 _06919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08694_ _01175_ _01178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_75_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13243__A1 _04255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09430__I _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09315_ _01730_ _01733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13794__A2 _05796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14991__A1 filters.filt_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09246_ _01676_ _01677_ _01669_ _01678_ _01679_ _01680_ _01681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_146_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09177_ channels.lfsr\[2\]\[5\] _01621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_32_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14743__A1 _06712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11557__A1 _03675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17564__CLK clknet_5_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_151_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_151_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11021__A3 _03243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15299__A2 _06955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput24 net24 bus_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_3_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11070_ filters.sample_filtered\[3\] _03291_ _03292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10021_ channels.atk_dec3\[6\] _02302_ _02303_ _02306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09922__A1 channels.sus_rel2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16799__A2 _01817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09605__I _01833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12809__A1 _04787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12031__I _04077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14760_ _06749_ _06733_ _06750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_11972_ _04044_ _04045_ _04046_ _04047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__13482__A1 _04480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13711_ _05712_ _05713_ _05714_ _05715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__10296__A1 _01307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10923_ channels.sample2\[11\] _03156_ _03161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14691_ _06515_ _06597_ _06686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_158_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16430_ _07818_ _08232_ _08233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_67_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13642_ filters.low\[1\] _05647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_175_3630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10854_ _03054_ _03104_ _03106_ _00279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_168_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_156_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09340__I _01013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10048__A1 _02324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16361_ channels.ch3_env\[3\] _08179_ _08183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13573_ _05461_ _05493_ _05578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__14982__A1 filters.high\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10785_ _03039_ _02939_ _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_136_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15312_ _07197_ _07201_ _07251_ _07270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_164_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_136_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12524_ _03333_ _04529_ _04522_ _04530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_16292_ _08143_ _00680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_171_3549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13797__I _04471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14734__A1 _06689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15243_ _07182_ _07186_ _07205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_152_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12455_ _04456_ _04460_ _04461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_124_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11406_ _01240_ _03582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_10_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15174_ _07135_ _07138_ _07139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_22_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12386_ _04258_ _04392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_50_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__16487__A1 _08274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14125_ _06123_ _06051_ _06124_ _06125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11337_ channels.adsr_state\[0\]\[1\] channels.adsr_state\[1\]\[1\] channels.adsr_state\[2\]\[1\]
+ channels.adsr_state\[3\]\[1\] _01147_ _01161_ _03531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_123_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14056_ _06022_ _06056_ _06057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11268_ filters.band\[15\] _03477_ _03236_ _03478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_123_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_37_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13007_ _05011_ _05012_ _05013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10219_ _01520_ _02478_ _02440_ _02479_ _02480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_27_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11199_ _03311_ _03379_ _03313_ _03412_ _03413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_94_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11720__B2 channels.atk_dec2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17746_ _00816_ clknet_leaf_55_clk tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14958_ _06928_ _06929_ _06921_ _06931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13473__A1 _03350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09141__A2 _01588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13909_ _04406_ _04929_ _05465_ _05466_ _05911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_89_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17677_ _00747_ clknet_leaf_61_clk tt_um_rejunity_sn76489.tone\[2\].gen.counter\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14889_ _06851_ _06867_ _06868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_134_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16628_ _01668_ _08386_ _08387_ _01670_ _00772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_175_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10039__A1 _02299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10396__I _02544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16559_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[2\] _08282_ _08339_ _08340_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09100_ _01547_ _01518_ _01552_ _01525_ _00075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_116_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09031_ _01479_ _01482_ _01490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11539__A1 _03662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_96_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10211__A1 channels.pw1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_57_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09933_ _02242_ _02235_ _02244_ _00220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_74_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_74_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09864_ _02185_ _02194_ _02197_ _00198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08815_ _01287_ _01288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09795_ _02112_ _02142_ _02147_ _00179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_29_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08746_ _01217_ _01227_ _01228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13464__A1 _05158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15590__C _06177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08677_ _01160_ _01161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_166_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15205__A2 _07168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09160__I _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_153_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10570_ _02790_ _02829_ _02830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_36_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_91_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09229_ channels.lfsr\[1\]\[11\] _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12240_ _04233_ _04245_ _04246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_131_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10202__A1 _01469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12171_ _03311_ _03312_ _03313_ filters.high\[6\] _04177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_0_31_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11950__A1 _04019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11122_ _03338_ _03340_ _03341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_120_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15930_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[2\] _07808_ _07812_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11053_ _03274_ _03275_ _03276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10004_ channels.atk_dec3\[0\] _02292_ _02294_ _02295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_73_Right_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15861_ _07724_ _07733_ spi_dac_i.counter\[4\] _07744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15781__B _07684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17600_ _00670_ clknet_leaf_40_clk spi_dac_i.spi_dat_buff_0\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14812_ _06778_ _06787_ _06734_ _06798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_157_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15792_ _07691_ _07692_ _00631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_153_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17531_ _00601_ clknet_leaf_82_clk filters.sample_buff\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_54_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11466__B1 _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14743_ _06712_ _06726_ _06734_ _06735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_11955_ _03866_ _04023_ _03862_ _04033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_58_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17462_ _00532_ clknet_leaf_2_clk filters.band\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10906_ channels.sample2\[4\] _03150_ _03151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08882__A1 channels.freq3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14674_ _04820_ _05370_ _06669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11886_ _03961_ _03971_ _03972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16413_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[10\] _08220_ _08221_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13625_ _04485_ _04884_ _05630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_17393_ _00463_ clknet_leaf_129_clk channels.env_counter\[2\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10837_ _03031_ _02890_ _03090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_15_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_82_Right_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_15_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16344_ _08172_ _00703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13556_ _05449_ _05561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14007__I0 filters.high\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10768_ _02992_ _02998_ _03023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12507_ _04512_ _04302_ _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16275_ _08129_ _08134_ _00672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_125_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13487_ _05475_ _05492_ _05493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_81_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10699_ _02501_ _02955_ _02956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15226_ _03411_ _07187_ _07189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12438_ _04443_ _04444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14860__B _06775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_247_clk clknet_5_0__leaf_clk clknet_leaf_247_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15157_ _07121_ _07097_ _05425_ _07122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_26_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12369_ _04374_ _04375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_121_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10744__A2 _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14108_ _06031_ _06032_ _06108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_91_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15088_ _04992_ _07012_ _07056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_91_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_91_Right_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14039_ _06037_ _06038_ _06039_ _06040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__13694__A1 _04694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input1_I addr[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09245__I _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08600_ channels.lfsr\[3\]\[4\] _01111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09580_ filters.mode_vol\[3\] _01790_ _01868_ channels.sus_rel2\[3\] _01968_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13446__A1 _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08531_ _01054_ _00003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_17729_ _00799_ clknet_leaf_60_clk tt_um_rejunity_sn76489.control_tone_freq\[2\]\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13997__A2 _05935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15710__I _07631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09014_ _01436_ _01473_ _01474_ _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_115_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_238_clk clknet_5_16__leaf_clk clknet_leaf_238_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_131_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13921__A2 _05208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09916_ _02216_ _02232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12488__A2 _04482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_8_clk_I clknet_5_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09847_ _02184_ _02185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_146_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09778_ channels.atk_dec1\[5\] _02134_ _02129_ _02136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09105__A2 _01556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08729_ _01199_ _01205_ _01206_ _01211_ _01213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_107_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16917__S _00987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_124_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11740_ _01150_ _03831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_124_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16926__A2 _00993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11671_ channels.sus_rel1\[4\] _01294_ _03762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_3_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13204__A4 _05145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13410_ _05405_ _05415_ _05416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_154_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10622_ channels.sample3\[2\] _02784_ _02881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14390_ _06372_ _06387_ _06388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_91_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13341_ _05259_ _05347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_84_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10553_ _02811_ _02812_ _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_51_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_180_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10974__A2 _03194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16060_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[1\] _07905_ _07939_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13272_ net48 _05276_ _05277_ _05278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_10484_ _02631_ _02639_ _02745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_leaf_229_clk clknet_5_17__leaf_clk clknet_leaf_229_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15011_ _04158_ _04776_ _06981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12223_ _04228_ _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__12715__A3 _04376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11923__A1 _02356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12154_ _04159_ _04160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_166_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15067__I _07030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11105_ _03321_ _03324_ _03325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_21_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12085_ _04056_ _04119_ _04123_ _00493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13676__A1 _05604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16962_ _00041_ clknet_leaf_233_clk channels.env_vol\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_34_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15913_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[3\] _07790_ _07795_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_159_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11036_ filters.sample_filtered\[1\] _03259_ _03260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11687__B1 _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16893_ _00957_ channels.exp_periods\[1\]\[0\] _00975_ _00976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15844_ _04776_ _07721_ _07730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15775_ _07295_ _07631_ _07648_ _07680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12987_ _04975_ _04989_ _04993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_14726_ _06718_ _06719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17514_ _00584_ clknet_leaf_21_clk filters.high\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11938_ _04001_ _04019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17445_ _00515_ clknet_leaf_147_clk channels.accum\[3\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10662__A1 _02402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14657_ _06613_ _06617_ _06651_ _06652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08950__S1 _01163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_25_Left_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__16626__I _08380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11869_ _03950_ _03951_ _03956_ _03750_ _03957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_172_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13608_ _04317_ _04713_ _05613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_157_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17376_ _00446_ clknet_leaf_207_clk channels.env_vol\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_172_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14588_ _04820_ _05280_ _06584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_31_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16327_ channels.env_vol\[1\]\[2\] _08160_ _08163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13539_ _05543_ _05544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16258_ filters.sample_buff\[7\] _08115_ _08122_ spi_dac_i.spi_dat_buff_0\[3\] spi_dac_i.spi_dat_buff_0\[4\]
+ _08119_ _08124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__14156__A2 _06155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15686__B _07573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12167__A1 filters.res_lut\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15209_ filters.high\[10\] _06934_ _07170_ _07172_ _07173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_113_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16189_ _08062_ _08043_ _08063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_34_Left_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15656__A2 _07579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16853__A1 _02707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09701_ _01777_ _02074_ _02080_ _00152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__16605__A1 _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09632_ _01995_ _02017_ _02018_ _00145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13419__A1 _05379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09563_ _01950_ _01951_ _01952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09099__A1 _01300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14092__A1 _04561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08514_ _01040_ _01030_ _00129_ _01041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09494_ _01884_ _01885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_43_Left_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12642__A2 _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15592__A1 channels.sample1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_144_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15344__A1 _07277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09023__A1 _01479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_52_Left_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_83_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_1300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11629__B _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_148_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10184__A3 channels.pw3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12705__I0 filters.high\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11133__A2 _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12910_ _04855_ _04856_ _04916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_6_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13890_ _05891_ _05892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_161_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12881__A2 _04332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12841_ _04220_ _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10892__A1 _02056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_61_Left_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15560_ _01932_ _07498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_167_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12772_ _04593_ _04777_ _04778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08837__A1 _01146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13830__A1 _05730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12633__A2 _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14511_ _03380_ _06080_ _06507_ _06187_ _00535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_11723_ _03813_ _03814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_16_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10644__A1 _02553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15491_ _06978_ _07435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_84_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13071__S _03185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17230_ _00300_ clknet_leaf_173_clk channels.sample1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_127_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14442_ _04355_ _05774_ _06439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_182_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11654_ _03131_ _03745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_181_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17161_ _00231_ clknet_leaf_121_clk channels.pw3\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10605_ _02858_ _02863_ _02864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_4_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14373_ _06347_ _06370_ _06371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11585_ _03640_ _01896_ _03695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_36_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16112_ _07988_ _07881_ _07989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10947__A2 _03104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13324_ _05329_ _05325_ _05330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_17092_ _00162_ clknet_leaf_110_clk channels.ctrl_reg1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_162_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10536_ _02747_ _02754_ _02796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_40_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15335__A1 filters.low\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_70_Left_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_165_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16043_ _07838_ _07920_ _07922_ _00652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09014__A1 _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13255_ _04185_ _05260_ _05261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_108_Right_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10467_ _02688_ _02690_ _02692_ _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12206_ _04206_ _04205_ _04211_ _04212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_126_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13186_ _05166_ _05191_ _05192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_10398_ _02656_ _02658_ _02659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10175__A3 channels.pw3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12214__I _04219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_214_clk_I clknet_5_21__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12137_ _04150_ _00518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13649__A1 _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12068_ _04103_ _04113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16945_ _00024_ clknet_leaf_227_clk channels.lfsr\[3\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12321__A1 _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11019_ _03241_ _03244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16876_ _00939_ _00962_ _00963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12872__A2 _04827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_229_clk_I clknet_5_17__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15827_ _03194_ _07628_ _07715_ _00643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_56_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08828__A1 channels.freq3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15758_ _03422_ _07633_ _07648_ _07668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_172_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_176_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08923__S1 _01162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14709_ _06700_ _06703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_15689_ filters.sample_filtered\[15\] _07602_ _07617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_172_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17428_ _00498_ clknet_leaf_159_clk channels.adsr_state\[2\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_145_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_109_Left_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_17359_ _00429_ clknet_leaf_172_clk channels.pw3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_60_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14129__A2 _05077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15326__A1 filters.low\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13888__A1 _04561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15629__A2 _07554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08994_ _01450_ _01447_ _01455_ _01456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_48_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_143_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_1197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12863__A2 _04844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09615_ channels.sus_rel2\[4\] _01936_ _02001_ channels.freq2\[4\] _02002_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11184__B _03398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_104_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15801__A2 _07697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09546_ channels.ctrl_reg3\[2\] _01882_ _01862_ channels.pw2\[10\] _01935_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_5_28__f_clk_I clknet_3_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09477_ _01832_ _01846_ _01868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_78_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09492__B2 channels.ctrl_reg3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15565__A1 channels.sample1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_164_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11370_ _03138_ _01333_ _03560_ _00341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_104_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10321_ _01157_ _02581_ _02582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11729__I1 channels.sus_rel1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13040_ _05014_ _05004_ _05045_ _05046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_10252_ _02512_ _02513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16817__A1 _01741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11354__A2 _01581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10183_ _02397_ _01098_ channels.pw2\[6\] _02444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_163_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_3721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_3732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14991_ filters.filt_2 filters.filt_1 channels.sample1\[2\] channels.sample2\[2\]
+ _06962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_16730_ tt_um_rejunity_sn76489.latch_control_reg\[1\] _08462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_13942_ _04186_ _05943_ _05944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16661_ _08333_ _08406_ _08407_ _08408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_13873_ _05846_ _05848_ _05875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_80_clk_I clknet_5_9__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15612_ _07486_ _07545_ _07546_ _07547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12824_ _04794_ _04795_ _04830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_69_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16592_ _08280_ _08362_ _08366_ _08367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_158_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13803__A1 _04221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15543_ filters.sample_buff\[2\] _07461_ _07451_ _07482_ _07483_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_178_3683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12755_ _04754_ _04757_ _04760_ _04761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_178_3694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11706_ _03795_ _03796_ _03785_ _03797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_56_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10093__A2 _02356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15474_ _06882_ _07415_ _07418_ _07419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__14359__A2 _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12686_ _04431_ _04519_ _04558_ _04690_ _04691_ _04692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA_clkbuf_leaf_95_clk_I clknet_5_13__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_139_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14425_ _04923_ _05732_ _06422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17213_ _00283_ clknet_leaf_170_clk channels.sample2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_182_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11637_ _03730_ _03731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13031__A2 _04992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17144_ _00214_ clknet_leaf_123_clk channels.sus_rel2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_141_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14356_ filters.band\[27\] _04578_ _06354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11568_ _03662_ _03680_ _03684_ _00415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_123_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13307_ _05307_ _05312_ _05313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_17075_ _00145_ clknet_leaf_119_clk net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10519_ _02763_ _02779_ _02780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_14287_ _06283_ _06285_ _06286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11499_ channels.freq1\[5\] _03633_ _03634_ _03636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16026_ _07814_ _07905_ _07906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09538__A2 _01904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13238_ _05178_ _05189_ _05243_ _05244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_122_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14531__A2 _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_153_clk_I clknet_5_29__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16808__A1 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[2\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13169_ _05069_ _04404_ _05175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_33_clk_I clknet_5_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16928_ tt_um_rejunity_sn76489.control_noise\[0\]\[1\] _00993_ _02272_ _00995_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_137_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_168_clk_I clknet_5_25__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12845__A2 _04850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09253__I _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_49_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_48_clk_I clknet_5_10__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16859_ _00944_ _00946_ _00947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_177_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09400_ _01757_ _01793_ _01797_ _00134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_137_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_94_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09331_ _01705_ _01736_ _01737_ _01708_ _00121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_73_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09474__A1 _01748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09474__B2 channels.pw2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13270__A2 _05188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13503__I _04848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11281__A1 filters.cutoff_lut\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_117_Left_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09262_ _01690_ _01683_ _01694_ _01674_ _00095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_30_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_62_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_157_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16814__I _00914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_106_clk_I clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09193_ channels.lfsr\[0\]\[6\] _01635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14334__I _04355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_141_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_1195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08977_ channels.freq3\[10\] _01439_ _01440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14286__A1 _03347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14038__A1 _05516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10102__I _02364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14589__A2 _05626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10870_ _03108_ _03121_ _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_116_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09529_ _01911_ _01912_ _01917_ _01918_ _01919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__11642__B _03735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08899__S0 _01146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12540_ _04172_ _04210_ _04533_ _04546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_176_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_156_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12471_ _04178_ _04477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_173_3591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14210_ _06207_ _06208_ _06209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_124_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11422_ _01103_ _03590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15190_ _07130_ _07131_ _07154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10378__A3 _02638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12772__A1 _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14141_ _06045_ _06053_ _06141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11353_ channels.ctrl_reg2\[0\] _01282_ _03547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_134_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09338__I _01740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10304_ _02548_ _02563_ _02565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14072_ _03472_ _06073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_11284_ net14 _03490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__15784__B _07684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12524__A1 _03333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13023_ _05024_ _05027_ _05029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_10235_ _01263_ _02495_ _02496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10166_ _01272_ _02427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12699__I _04476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17762_ _00832_ clknet_5_9__leaf_clk tt_um_rejunity_sn76489.clk_counter\[0\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14974_ _06922_ _06945_ _06946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_10097_ _02360_ _01569_ _02361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16713_ _02100_ _08450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13925_ _05922_ _05926_ _05927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_17693_ _00763_ clknet_leaf_217_clk channels.lfsr\[0\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16644_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[9\] tt_um_rejunity_sn76489.tone\[0\].gen.counter\[8\]
+ _08391_ _08392_ _08393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_13856_ _05757_ _05858_ _05859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_159_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12807_ _04799_ _04808_ _04809_ _04813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_16575_ _08349_ _08352_ _08353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_29_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13787_ _04966_ _04447_ _05622_ _05790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_44_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10999_ _03223_ _03224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_139_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12738_ _04738_ _04741_ _04743_ _04744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_15526_ channels.sample1\[1\] _03335_ _07467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11802__A3 _03887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15457_ _07402_ _07403_ _00585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12669_ _04610_ _04627_ _04675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__11015__A1 filters.hp vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14408_ _06373_ _06386_ _06405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11015__B2 filters.bp vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_160_Right_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15388_ _07324_ _07338_ _07339_ _07340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__14752__A2 _06731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17127_ _00197_ clknet_leaf_127_clk channels.ctrl_reg2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14339_ _06335_ _06213_ _06336_ _06337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__10682__I _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17058_ _00128_ clknet_leaf_76_clk filters.res_filt\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14504__A2 _03378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16009_ _07884_ _07888_ _07889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08900_ _01367_ _01368_ _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09880_ _02160_ _02201_ _02207_ _00204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_148_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08831_ _01188_ _01304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_100_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08762_ _01240_ _01241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08693_ channels.exp_periods\[0\]\[0\] channels.exp_periods\[1\]\[0\] _01176_ _01177_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08498__A2 _01019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13491__A2 _05354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_137_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13243__A2 _04392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09314_ _01728_ _01732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_119_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12597__A4 _04601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14991__A2 filters.filt_1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09245_ _01606_ _01680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_91_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09176_ _01616_ _01611_ _01620_ _01599_ _00083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_133_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12754__A1 _04641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_151_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_151_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09158__I _01604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput25 net25 bus_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_112_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10020_ _02238_ _02301_ _02305_ _00246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__14259__A1 _06142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11971_ _03914_ _04039_ _04046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_98_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13482__A2 _05487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13710_ _04449_ _04945_ _05714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13344__S _04710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11493__A1 _03515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10922_ _02365_ _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14690_ _06653_ _06662_ _06684_ _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__15759__A1 _06714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_158_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13641_ _05644_ _05645_ _05646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_116_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10853_ channels.sample3\[8\] _03105_ _03106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13234__A2 _05234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_175_3631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16360_ _03954_ _08177_ _08182_ _00709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13572_ _05565_ _05576_ _05577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10784_ _02676_ _03039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_67_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14982__A2 _06934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15311_ _03467_ _06910_ _07268_ _07269_ _00573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_136_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12993__A1 _04211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12523_ _04175_ _04529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16291_ channels.env_counter\[3\]\[1\] _08143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__16454__I _07683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15242_ _07182_ _07186_ _07204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12454_ _04457_ _04458_ _04459_ _04460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_48_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_1168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11405_ _01089_ _03581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_62_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15173_ _07098_ _07136_ _07137_ _07138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_10_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12385_ _04388_ _04390_ _04391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_151_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09068__I _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14124_ _06049_ _06050_ _06124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_104_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11336_ _03529_ _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10220__A2 _02473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14055_ _06024_ _06055_ _06056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_11267_ _03476_ _03477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13006_ _04984_ _04983_ _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_37_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10218_ channels.pw1\[4\] _02435_ _02479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_37_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11198_ filters.band\[11\] _03412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_20_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12222__I _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10149_ _02397_ _01250_ channels.pw2\[8\] _02410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_27_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17745_ _00815_ clknet_leaf_55_clk tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09677__A1 channels.freq1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14957_ _06921_ _06928_ _06929_ _06930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09677__B2 channels.sus_rel2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13473__A2 _04192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13908_ _04406_ _05909_ _05466_ _04929_ _05910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_17676_ _00746_ clknet_leaf_80_clk tt_um_rejunity_sn76489.tone\[2\].gen.counter\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14888_ _06864_ _06866_ _06867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_43_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16627_ _08382_ _08387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09429__A1 _01819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13839_ _05827_ _05841_ _05842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_119_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16558_ _01752_ _08339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_70_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13988__I _05796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15509_ _07450_ _07451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_150_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16489_ _08280_ _08281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09030_ channels.accum\[0\]\[14\] _01489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_155_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16478__A2 _08267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09932_ channels.sus_rel2\[7\] _02236_ _02243_ _02244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_74_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13161__A1 _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09863_ channels.ctrl_reg2\[1\] _02195_ _02189_ _02197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08814_ _01286_ _01287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09794_ channels.sus_rel1\[2\] _02143_ _02146_ _02147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08745_ _01186_ _01222_ _01227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13464__A2 _05469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11475__A1 _03612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08676_ _01159_ _01160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_95_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14413__A1 _06314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08891__A2 _01360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11920__B _01585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_153_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09228_ channels.lfsr\[0\]\[11\] _01665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_106_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09159_ _01304_ _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_131_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11211__I _03395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12170_ _04175_ _04176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_11121_ _03321_ _03324_ _03339_ _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_102_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15141__A2 channels.sample2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11052_ filters.high\[2\] _03209_ _03275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10003_ _02293_ _02294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15860_ _07742_ _07743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_129_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14811_ _06779_ _06796_ _06788_ _06797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_15791_ _07327_ _07682_ _07684_ _07692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09659__B2 channels.ctrl_reg3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14652__A1 filters.band\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17530_ _00600_ clknet_leaf_82_clk filters.sample_buff\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11954_ _03862_ _03866_ _04023_ _04032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_118_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_98_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14742_ _06716_ _06734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_93_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10905_ _03149_ _03150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_169_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14673_ _04806_ _05663_ _06668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17461_ _00531_ clknet_leaf_1_clk filters.band\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11885_ _03541_ _03752_ _03971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xclkbuf_leaf_192_clk clknet_5_23__leaf_clk clknet_leaf_192_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_156_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16412_ _08197_ _08220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_156_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13624_ _05485_ _05627_ _05628_ _05629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10836_ _03088_ _02840_ _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17392_ _00462_ clknet_leaf_130_clk channels.env_counter\[2\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14955__A2 _06912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13555_ _04645_ _05560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_16343_ _01225_ _01255_ _01258_ channels.exp_counter\[0\]\[1\] _08172_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10767_ _03000_ _03003_ _03022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_82_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09831__A1 channels.freq2\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14007__I1 filters.band\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12506_ _04511_ _04512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_81_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16274_ filters.sample_buff\[13\] _07742_ _08130_ spi_dac_i.spi_dat_buff_0\[9\] spi_dac_i.spi_dat_buff_0\[10\]
+ _08096_ _08134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_13486_ _05477_ _05491_ _05492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10698_ _02576_ _02955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_124_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12718__A1 _04458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15225_ filters.low\[11\] _07187_ _07188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_12437_ filters.cutoff_lut\[11\] _04442_ _04443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_125_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09595__B1 _01954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15156_ _05379_ _05403_ _07121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12368_ filters.cutoff_lut\[10\] filters.res_lut\[10\] _04166_ _04374_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14107_ _06036_ _06040_ _06106_ _06107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11319_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[3\] _03509_ _03517_ _03518_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_121_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10960__I _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15087_ _07052_ _07054_ _07055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_91_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12299_ _04289_ _04304_ _04305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_129_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13143__A1 _04278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14038_ _05516_ _05230_ _06039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09898__A1 channels.atk_dec2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13694__A2 _05075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14891__A1 _06520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13048__I _04946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_173_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12887__I _04316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15989_ _07869_ _07870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_136_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08530_ _01047_ _01053_ _01054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_17728_ _00798_ clknet_leaf_60_clk tt_um_rejunity_sn76489.control_tone_freq\[2\]\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17659_ _00729_ clknet_leaf_49_clk tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14808__S _03472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_98_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10283__I2 channels.ch3_env\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09013_ _01465_ _01457_ _01472_ _01474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__12709__A1 _04274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10196__A1 channels.pw1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09915_ _02188_ _02227_ _02231_ _00215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09889__A1 channels.atk_dec2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13685__A2 _05260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09846_ _01755_ _02184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11696__A1 _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_146_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09777_ _01801_ _02133_ _02135_ _00173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_154_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12797__I _04783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14634__A1 _04447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08728_ _01199_ _01205_ _01206_ _01211_ _01212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_90_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11448__A1 _03600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_124_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08659_ _01142_ _01143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_87_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10120__A1 channels.ctrl_reg3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_174_clk clknet_5_24__leaf_clk clknet_leaf_174_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_139_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10120__B2 channels.ctrl_reg2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11670_ _03748_ _03759_ _03760_ _03761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_3_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10621_ _02835_ _02879_ _02880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_113_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09813__A1 channels.sus_rel1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_12_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13340_ _05341_ _05345_ _05346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_36_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08515__I net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11620__A1 _03666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10552_ _02535_ _02500_ _02812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13271_ _05184_ _05188_ _05277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__16732__I _08463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10483_ _02742_ _02649_ _02743_ _02744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_121_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15010_ filters.high\[4\] _06955_ _06980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09577__B1 _01964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12222_ _04227_ _04228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_60_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12153_ _04158_ _03226_ _04159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__09346__I _01013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11104_ _03322_ _03307_ _03323_ _03324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_12084_ channels.env_counter\[0\]\[10\] _04120_ _04123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16961_ _00040_ clknet_leaf_213_clk channels.env_vol\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_34_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15912_ _07793_ _07794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_95_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11035_ _03257_ _03258_ _03259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_159_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16892_ _00974_ _00975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11687__B2 _03777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08552__A1 _01062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15843_ _07718_ _07729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_99_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12986_ _04952_ _04991_ _04992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_15774_ _07678_ _07679_ _00626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_24_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17513_ _00583_ clknet_leaf_21_clk filters.high\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14725_ _06717_ _06718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_11937_ _04008_ _04017_ _04018_ _00450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_165_clk clknet_5_25__leaf_clk clknet_leaf_165_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17444_ _00514_ clknet_leaf_151_clk channels.accum\[3\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14656_ _06618_ _06636_ _06650_ _06651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_11868_ _03536_ _03951_ _03956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13607_ _04377_ _04751_ _05612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10819_ _03061_ _03072_ _03073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_83_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17375_ _00445_ clknet_leaf_204_clk channels.env_vol\[0\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_156_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11799_ _03835_ _03890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_144_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14587_ _06581_ _06423_ _06582_ _06583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_43_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16326_ _03948_ _08158_ _08162_ _00695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13538_ _03730_ _03477_ _05543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_31_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16257_ _08121_ _08123_ _00665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13469_ _05474_ _05464_ _05475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_93_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09568__B1 _01866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15208_ _06909_ _07171_ _07172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16188_ _08017_ _08021_ _08062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_26_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15139_ _07102_ _07103_ _07104_ _07105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__13116__A1 _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09700_ channels.freq1\[11\] _02075_ _02077_ _02080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_156_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11678__A1 channels.sus_rel3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09631_ _01934_ net26 _01809_ _02018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16605__A2 _08374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13419__A2 _05403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09562_ channels.ctrl_reg2\[2\] _01829_ _01879_ channels.freq2\[2\] _01951_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_69_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08513_ _01008_ _01040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09493_ _01854_ _01860_ _01884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_136_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16369__A1 channels.ch3_env\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_156_clk clknet_5_29__leaf_clk clknet_leaf_156_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_33_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11850__A1 _03744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_102_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11602__A1 channels.pw3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12650__I0 _04644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09023__A2 _01482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14072__I _03472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08782__A1 _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12705__I1 filters.band\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12330__A2 _04219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09829_ channels.freq2\[12\] _02171_ _02167_ _02172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_126_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12881__A3 _04800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12840_ _04790_ _04797_ _04845_ _04846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_17_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12771_ filters.cutoff_lut\[11\] _04776_ _04777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12094__A1 _01240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_147_clk clknet_5_29__leaf_clk clknet_leaf_147_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_55_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11722_ _03533_ _03808_ _03810_ _03812_ _03813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_14510_ _06403_ _06506_ _06507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_15490_ _07426_ _07432_ _07433_ _07434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10644__A2 _02575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11653_ _01319_ _03744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_126_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14441_ _06436_ _06328_ _06437_ _06438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_138_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13594__A1 _05594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10604_ _02859_ _02862_ _02863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_17160_ _00230_ clknet_leaf_166_clk channels.pw3\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14372_ _06350_ _06369_ _06370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11584_ _03677_ _03687_ _03694_ _00421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_65_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15787__B _07684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09262__A2 _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16111_ _07795_ _07988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13323_ _05326_ _05327_ _05328_ _05329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_51_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10535_ _02747_ _02754_ _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_36_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17091_ _00161_ clknet_leaf_110_clk channels.ctrl_reg1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_52_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13346__A1 _04184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16042_ spi_dac_i.spi_dat_buff_1\[1\] _07867_ _07921_ spi_dac_i.spi_dat_buff_1\[2\]
+ _07871_ _07922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_13254_ _05259_ _05260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_161_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10466_ _02696_ _02702_ _02719_ _02726_ _02727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_122_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12205_ _04208_ _04211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_86_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13185_ _05168_ _05171_ _05190_ _05191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_62_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10397_ _02655_ _02657_ _02569_ _02658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_12136_ channels.accum\[3\]\[16\] _04150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10015__I _02290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12067_ _04025_ _04105_ _04112_ _00486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16944_ _00023_ clknet_leaf_227_clk channels.lfsr\[3\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11018_ _03242_ _03243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12321__A2 _04326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16599__A1 _08356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16875_ _01211_ _00955_ _00961_ _00962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_95_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12230__I _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15826_ _03735_ _07714_ _07715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_138_clk clknet_5_31__leaf_clk clknet_leaf_138_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15757_ _06695_ _07632_ _07667_ _00621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_12969_ _04961_ _04964_ _04974_ _04975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_14708_ _06701_ _06691_ _06702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_47_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15688_ filters.sample_buff\[13\] _03452_ _07602_ _07616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_47_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17427_ _00497_ clknet_leaf_129_clk channels.env_counter\[0\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_142_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14639_ _06629_ _06630_ _06633_ _06634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_64_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17358_ _00428_ clknet_leaf_95_clk channels.pw3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16309_ channels.env_counter\[3\]\[10\] _08152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_126_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_60_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17289_ _00359_ clknet_leaf_161_clk channels.accum\[2\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08993_ _01453_ _01454_ _01455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_103_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16321__B _01821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15716__I _07636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_143_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09614_ _01880_ _02001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_104_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15262__A1 filters.high\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_104_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09545_ _01874_ _01934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_129_clk clknet_5_30__leaf_clk clknet_leaf_129_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_167_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13812__A2 _05714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_174_Right_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09476_ _01866_ _01867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_4_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16762__A1 _01800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_119_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10320_ channels.env_vol\[0\]\[5\] channels.env_vol\[1\]\[5\] _02519_ _02581_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10251_ _02372_ _02510_ _02511_ _02512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_10182_ _02438_ _02442_ _02443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_163_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10562__A1 _01556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_180_3722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14990_ _06942_ _06960_ _06940_ _06961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_180_3733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09624__I _01954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13500__A1 _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13941_ filters.high\[24\] filters.band\[24\] _05179_ _05943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_156_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16660_ _08394_ _08405_ _08404_ _08407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13872_ _05846_ _05848_ _05874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15611_ _07537_ _07532_ _07544_ _07546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_12823_ _04794_ _04795_ _04829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_16591_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[8\] _08329_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[8\]
+ _08366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13803__A2 _05187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_141_Right_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15542_ _07480_ _07481_ _07482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_178_3684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12754_ _04641_ _04759_ _04760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_178_3695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11705_ channels.sus_rel3\[1\] _01077_ _01425_ channels.sus_rel2\[1\] _03796_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_127_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15473_ _07415_ _07417_ _07418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_12685_ _04556_ _04557_ _04691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_167_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17212_ _00282_ clknet_leaf_171_clk channels.sample3\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_139_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11636_ _03729_ _03730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_14424_ _05183_ _06027_ _06421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17143_ _00213_ clknet_leaf_128_clk channels.sus_rel2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_11567_ channels.freq3\[1\] _03681_ _03682_ _03684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14355_ _06351_ _06352_ _06353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10518_ _02767_ _02778_ _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13306_ _05308_ _05311_ _05312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_80_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17074_ _00144_ clknet_leaf_119_clk net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14286_ _03347_ _06177_ _06284_ _06285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_11498_ _02319_ _03632_ _03635_ _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_52_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16025_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[0\] _07809_ _07905_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_123_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13237_ _05172_ _05242_ _05177_ _05243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10449_ _02642_ _02710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13334__A4 _04712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13168_ _04228_ _04737_ _05174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12119_ _04141_ _00509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13099_ _03252_ _04224_ _04880_ _05105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_88_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16927_ _01741_ _00993_ _00994_ _00857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_137_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16858_ _03768_ _03747_ _00942_ _00945_ _00946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_15809_ _07383_ _07694_ _07695_ _07705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_137_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16789_ _03499_ _00897_ _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09330_ _01577_ _01736_ _01737_ _01703_ _00120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_172_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10608__A2 _02823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09474__A2 _01844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09261_ _01691_ _01692_ _01682_ _01693_ _01679_ _01680_ _01694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_62_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_62_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09192_ _01610_ _01634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_90_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09226__A2 _01659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11033__A2 _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08985__A1 _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13730__A1 _05730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08976_ _01397_ _01439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14286__A2 _06177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17638__CLK clknet_5_19__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15235__A1 _07146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09528_ channels.atk_dec3\[1\] _01867_ _01869_ channels.sus_rel2\[1\] _01871_ channels.freq3\[1\]
+ _01918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_79_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09465__A2 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08899__S1 _01161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09459_ net2 _01787_ _01850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16735__A1 _03710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_213_clk_I clknet_5_21__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_156_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13549__A1 _05444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_156_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12470_ _04227_ _04476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_152_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16226__B _08098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_3592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11421_ channels.accum\[1\]\[0\] _03589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_151_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12221__A1 filters.res_lut\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14140_ _06052_ _06140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_85_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11352_ _03534_ _03544_ _03546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_134_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_134_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_228_clk_I clknet_5_17__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10303_ _02548_ _02563_ _02564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14071_ _06070_ _06071_ _06072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11283_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[0\] _03489_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_131_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13022_ _05024_ _05027_ _05028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10234_ _01266_ channels.ctrl_reg2\[6\] _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12524__A2 _04529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10165_ _01249_ _02426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09354__I _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17761_ _00831_ clknet_leaf_70_clk tt_um_rejunity_sn76489.latch_control_reg\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14973_ _06922_ _06923_ _06925_ _06945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_10096_ _01085_ _02360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_89_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16712_ _01755_ _08449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13924_ _05923_ _05924_ _05925_ _05926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_17692_ _00762_ clknet_leaf_216_clk channels.lfsr\[0\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15226__A1 _03411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08900__A1 _01367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16643_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[7\] tt_um_rejunity_sn76489.tone\[0\].gen.counter\[6\]
+ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[5\] tt_um_rejunity_sn76489.tone\[0\].gen.counter\[4\]
+ _08392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_53_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13855_ _05548_ _05650_ _05858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12806_ _04746_ _04719_ _04812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_16574_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[5\] _08328_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[5\]
+ _08352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_97_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13786_ _05693_ _05787_ _05788_ _05789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_10998_ _03222_ _03223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_44_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15525_ channels.sample2\[1\] _03219_ _07465_ _03229_ _07466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_128_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12737_ _04510_ _04742_ _04743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12460__A1 _04319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15456_ filters.high\[27\] _06983_ _07333_ _07403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_84_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_155_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12668_ _04610_ _04627_ _04662_ _04673_ _04674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_26_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14407_ _06376_ _06385_ _06404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10963__I _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11015__A2 _03236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11619_ channels.pw2\[3\] _03713_ _03714_ _03718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15387_ _07328_ _07337_ _07339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12599_ _04261_ _04541_ _04605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_170_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17126_ _00196_ clknet_leaf_113_clk channels.pw2\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_13_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14338_ _06211_ _06212_ _06336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_151_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17057_ _00127_ clknet_leaf_89_clk filters.filt_3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14269_ _06265_ _06266_ _06268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16008_ _07885_ _07887_ _07888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_59_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08830_ _01301_ _01302_ _01303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_100_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08761_ _01083_ _01240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_164_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08692_ _01175_ _01176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_75_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_135_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09313_ _01638_ _01729_ _01731_ _01641_ _00109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12451__A1 _04366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14991__A3 channels.sample1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_60_clk clknet_5_8__leaf_clk clknet_leaf_60_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_145_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09244_ _01604_ _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_75_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_146_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11969__I _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09175_ _01617_ _01618_ _01609_ _01619_ _01605_ _01607_ _01620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_111_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13951__A1 _04392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_79_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_101_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput26 net26 bus_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_141_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_112_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14080__I _05544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_94_clk_I clknet_5_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08959_ _01414_ _01415_ _01423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11970_ _03914_ _04039_ _04045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15208__A1 _06909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10921_ _03154_ _03136_ _03159_ _00293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15759__A2 _07632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_158_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13640_ _05549_ _05550_ _05643_ _05645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10852_ _02974_ _03105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_5_12__f_clk_I clknet_3_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_3632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_152_clk_I clknet_5_29__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13571_ _05568_ _05575_ _05576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10783_ _02961_ _02873_ _03038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_51_clk clknet_5_10__leaf_clk clknet_leaf_51_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10453__B1 _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15310_ _06186_ _07269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_leaf_32_clk_I clknet_5_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12993__A2 _04966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12522_ _04521_ _04527_ _04528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_16290_ _08142_ _00679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_136_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15241_ _07202_ _07203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_109_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12453_ _03273_ _04372_ _04243_ _04459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__14255__I _05560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09349__I _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13942__A1 _04186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11404_ channels.accum\[2\]\[16\] _03580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_105_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12384_ _04389_ _04390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15172_ _03360_ _07111_ _07137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_151_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_136_Left_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_47_clk_I clknet_5_10__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14123_ _06049_ _06050_ _06123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11335_ channels.adsr_state\[0\]\[0\] channels.adsr_state\[1\]\[0\] channels.adsr_state\[2\]\[0\]
+ channels.adsr_state\[3\]\[0\] _01146_ _01160_ _03529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_123_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14498__A2 _06394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11266_ _03475_ _03476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_14054_ _06042_ _06054_ _06055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__10508__A1 _01542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09374__A1 _01767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13005_ _05008_ _05009_ _05010_ _05011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_94_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10217_ _01265_ _01098_ channels.pw2\[4\] _02478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_37_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11197_ filters.low\[11\] _03411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_20_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10148_ _02406_ _02407_ _02408_ _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_clkbuf_leaf_105_clk_I clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17744_ _00814_ clknet_leaf_54_clk tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10079_ _02328_ _02340_ _02346_ _00264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14956_ _05534_ _06915_ _06926_ _06929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_145_Left_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09812__I _01818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13473__A3 _05220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13907_ _05229_ _05909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17675_ _00745_ clknet_leaf_81_clk tt_um_rejunity_sn76489.tone\[2\].gen.counter\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14887_ _06854_ _06857_ _06865_ _06866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_58_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08980__S0 _01149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16626_ _08380_ _08386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_134_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13838_ _05832_ _05840_ _05841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_130_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16557_ _08333_ _08336_ _08337_ _08338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_13769_ _05770_ _05771_ _05772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_84_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_42_clk clknet_5_3__leaf_clk clknet_leaf_42_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_57_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15508_ _07449_ _07450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16488_ _08241_ _08280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_155_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15439_ _07372_ _07375_ _07374_ _07387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_154_Left_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_96_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17109_ _00179_ clknet_leaf_114_clk channels.sus_rel1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09931_ _02216_ _02243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_180_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_74_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09862_ _02179_ _02194_ _02196_ _00197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_141_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08813_ _01285_ _01286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_175_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09793_ _02137_ _02146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_163_Left_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09117__A1 _01300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15724__I _07332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08744_ _01226_ _00045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08675_ _01158_ _01159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_178_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12672__A1 _04674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_178_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14413__A2 _06346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_33_clk clknet_5_2__leaf_clk clknet_leaf_33_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_36_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_172_Left_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_134_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09227_ channels.lfsr\[2\]\[12\] _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_90_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_170_3540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_114_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09158_ _01604_ _01605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_131_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09089_ _01542_ _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__15677__A1 filters.sample_buff\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11120_ _03318_ _03319_ _03309_ _03339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_102_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11051_ _03268_ _03188_ _03273_ _03206_ _03274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_101_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_181_Left_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__15429__A1 _07373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10002_ _02174_ _02293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10910__A1 channels.sample2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_129_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14810_ _06757_ _06773_ _06796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15790_ _06809_ _07690_ _07691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09659__A2 _01871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14741_ _06713_ _06727_ _06733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11953_ _04027_ _04029_ _04031_ _00453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16929__A1 _08449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11466__A2 _01230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17460_ _00530_ clknet_leaf_249_clk filters.band\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10904_ _01103_ _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_157_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14672_ _06576_ _06665_ _06666_ _06589_ _06574_ _06667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_54_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11884_ _03540_ _03969_ _03970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16411_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[9\] _08212_ _08219_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_157_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13623_ _04473_ _05231_ _05624_ _05626_ _05628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_17391_ _00461_ clknet_leaf_123_clk channels.env_counter\[2\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10835_ _02994_ _03088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_94_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16342_ _08171_ _00702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13554_ _05459_ _05556_ _05557_ _05558_ _05456_ _05559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_137_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10766_ _03001_ _03002_ _03021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_66_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12505_ _04510_ _04511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_164_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16273_ _08129_ _08133_ _00671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_89_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13485_ _05482_ _05490_ _05491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10697_ _02555_ _02638_ _02954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09079__I _01533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12718__A2 _04459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15224_ _07179_ _07182_ _07186_ _07187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_164_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12436_ _04441_ _04442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_22_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09595__A1 filters.cutoff_lut\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09595__B2 channels.freq1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15155_ _03359_ _07064_ _07120_ _07089_ _00566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_164_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12367_ _04372_ _04321_ _04373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14106_ _06030_ _06035_ _06106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11318_ _03516_ _03517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_12298_ _04300_ _04303_ _04304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_15086_ _07053_ _05421_ _07054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_91_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14340__A1 _04326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13143__A2 _04780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14037_ _05469_ _04825_ _06038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11249_ _03236_ _03458_ _03459_ _03460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__10181__C _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15988_ _07868_ _07869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_179_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17727_ _00797_ clknet_leaf_60_clk tt_um_rejunity_sn76489.control_tone_freq\[2\]\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14939_ _06908_ _06913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_77_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17658_ _00728_ clknet_leaf_51_clk tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15199__A3 _07162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16609_ _01598_ _08376_ _08379_ _01601_ _00761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_17589_ _00659_ clknet_leaf_44_clk spi_dac_i.spi_dat_buff_1\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_15_clk clknet_5_6__leaf_clk clknet_leaf_15_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_161_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09012_ _01465_ _01457_ _01472_ _01473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_116_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12709__A2 _04295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15719__I _07639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15659__A1 channels.sample2\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09914_ channels.sus_rel2\[2\] _02228_ _02224_ _02231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10091__C _02354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09845_ _02179_ _02181_ _02183_ _00193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_146_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09776_ channels.atk_dec1\[4\] _02134_ _02129_ _02135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08727_ _01174_ _01207_ _01210_ _01211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_107_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_107_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08658_ _01141_ _01142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_87_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08589_ _01104_ _01105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10620_ _02837_ _02878_ _02879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_92_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10551_ _02544_ _02554_ _02811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12318__I _04323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10482_ _02627_ _02640_ _02743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13270_ _05184_ _05188_ _05276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09577__A1 channels.sus_rel3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14570__A1 _04446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12221_ filters.res_lut\[5\] _04167_ _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_4
XANTENNA__09577__B2 channels.sus_rel1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12152_ _01093_ _04158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_11103_ filters.sample_filtered\[4\] _03304_ _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14322__A1 _05469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12083_ _04051_ _04119_ _04122_ _00492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16960_ _00039_ clknet_leaf_211_clk channels.env_vol\[3\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15911_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[0\] _07790_ _07793_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_34_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11034_ filters.high\[1\] _03209_ _03258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16891_ _01724_ _00973_ _00974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__11687__A2 _03755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15842_ _07727_ _07728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15773_ filters.low\[16\] _07670_ _07671_ _07679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12985_ _04975_ _04989_ _04990_ _04991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__12002__B _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17512_ _00582_ clknet_leaf_27_clk filters.high\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_169_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10301__I _02561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08935__S0 _01148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14724_ _06716_ _06717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_11936_ channels.env_counter\[2\]\[1\] _04013_ _04018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17443_ _00513_ clknet_leaf_146_clk channels.accum\[3\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14389__A1 _06373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14655_ _06639_ _06649_ _06650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11867_ _03939_ _03954_ _03955_ _00443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15050__A2 channels.sample2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13606_ _05158_ _05516_ _05611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13061__A1 _04705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17374_ _00444_ clknet_leaf_207_clk channels.env_vol\[0\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10818_ _03062_ _03071_ _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_14586_ _06421_ _06422_ _06582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_11798_ _03884_ _03885_ _03888_ _03889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16325_ channels.env_vol\[1\]\[1\] _08160_ _08162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_171_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13537_ _04161_ _05539_ _05542_ _00526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10414__A3 _02662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10749_ _02999_ _03004_ _03005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_131_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16256_ filters.sample_buff\[6\] _08115_ _08122_ spi_dac_i.spi_dat_buff_0\[2\] spi_dac_i.spi_dat_buff_0\[3\]
+ _08119_ _08123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_36_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13468_ _05468_ _05473_ _05474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_152_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09568__A1 filters.cutoff_lut\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15207_ _07169_ _07146_ _07149_ _07171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09568__B2 channels.atk_dec3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12419_ _04423_ _04424_ _04425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_16187_ _07997_ _08060_ _08046_ _07994_ _08061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_23_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13399_ _05391_ _05401_ _05405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_15138_ _07074_ _07075_ _07104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_121_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16798__C _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15069_ _07026_ _07036_ _07037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_4_clk clknet_5_4__leaf_clk clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_103_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_155_Right_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09630_ _02006_ _02016_ _02017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_136_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09561_ channels.pw1\[2\] _01884_ _01892_ channels.freq2\[10\] _01950_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11307__I _03507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08512_ _01039_ _00000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_19_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09492_ channels.freq2\[0\] _01880_ _01882_ channels.ctrl_reg3\[0\] _01883_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_176_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15041__A2 _06996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09256__B1 _01689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_5_18__f_clk clknet_3_4_0_clk clknet_5_18__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_2_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09103__S0 _01139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_148_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14304__A1 _06281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08782__A2 _01253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14304__B2 _06173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_165_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11669__A2 _03759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_109_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09828_ _02162_ _02171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_126_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_122_Right_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_126_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09182__I _01588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_161_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09759_ _01819_ _02116_ _02122_ _00168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10121__I _02381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12770_ _04442_ _04776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_output26_I net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11721_ _03791_ _03811_ _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14440_ _06326_ _06327_ _06437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_166_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11652_ _03742_ _03743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_182_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10603_ _02860_ _02861_ _02862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_64_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14371_ _06353_ _06368_ _06369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_153_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11583_ channels.freq3\[7\] _03688_ _03690_ _03694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_24_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16110_ _07824_ _07986_ _07987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13322_ _04315_ _04404_ _05328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17090_ _00160_ clknet_leaf_113_clk channels.pw1\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10534_ _02763_ _02779_ _02793_ _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_150_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16041_ _07868_ _07921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_134_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10465_ _02722_ _02723_ _02724_ _02725_ _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_13253_ filters.high\[18\] filters.band\[18\] _03185_ _05259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_161_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12204_ _04205_ _04209_ _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_110_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13184_ _05178_ _05189_ _05190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10396_ _02544_ _02657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_20_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12135_ _04149_ _00517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_159_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16943_ _00022_ clknet_leaf_226_clk channels.lfsr\[3\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12066_ channels.env_counter\[0\]\[3\] _04108_ _04112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12857__A1 _04400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15308__B _07086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09722__A1 _01757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11017_ _03214_ _03216_ _03241_ _03242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_16874_ _00946_ _00960_ _00940_ _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10332__A2 _02535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15825_ _03214_ _03216_ _03731_ _07714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_56_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15756_ _03411_ _07633_ _07648_ _07667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12968_ _04972_ _04973_ _04974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_157_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14707_ _06700_ _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_11919_ _01185_ _01191_ _01198_ _01223_ _04002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_158_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15687_ filters.sample_buff\[14\] _07615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_47_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12899_ _04901_ _04904_ _04905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_47_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17426_ _00496_ clknet_leaf_136_clk channels.env_counter\[0\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14638_ _06584_ _06631_ _06632_ _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_129_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17357_ _00427_ clknet_leaf_101_clk channels.pw3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_71_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14569_ _06440_ _06441_ _06564_ _06565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_83_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_172_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11596__A1 _03666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16308_ _08151_ _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17288_ _00358_ clknet_leaf_157_clk channels.accum\[2\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11797__I _03887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16239_ _08109_ _08110_ _00660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13337__A2 _04711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09267__I _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10020__A1 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09961__A1 _01781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08992_ channels.accum\[0\]\[11\] channels.accum\[1\]\[11\] channels.accum\[2\]\[11\]
+ channels.accum\[3\]\[11\] _01149_ _01165_ _01454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_76_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_103_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_76_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_143_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10323__A2 _02543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09613_ channels.freq3\[4\] _01937_ _01999_ channels.ctrl_reg3\[4\] _02000_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15262__A2 _07062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09544_ _01932_ _01933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_167_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09730__I _02101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_84_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09475_ _01825_ _01840_ _01866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_65_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14792__B _06765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13576__A2 _05520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_119_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13328__A2 _05263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14525__A1 _06520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10250_ _01508_ _02381_ _02511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08755__A2 _01230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10181_ _02439_ _01286_ _02440_ _02441_ _01520_ _02442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_163_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12839__A1 _04792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_180_3723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09704__A1 channels.freq1\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13940_ _04294_ _05504_ _05942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11511__A1 channels.pw1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13871_ _05743_ _05746_ _05873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__16738__I _08463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15610_ _07537_ _07532_ _07544_ _07545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_12822_ _04821_ _04827_ _04828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_69_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16590_ _08364_ _08365_ _00756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_97_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10078__A1 filters.cutoff_lut\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15541_ _07472_ _07473_ _07479_ _07481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_69_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12753_ _04758_ _04759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_69_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_3685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_178_3696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11704_ channels.atk_dec3\[1\] _01077_ _01425_ channels.atk_dec2\[1\] _03795_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_139_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15472_ _07416_ _06717_ _07417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_38_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12684_ _04684_ _04688_ _04689_ _04690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_37_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17211_ _00281_ clknet_leaf_94_clk channels.sample3\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_139_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14423_ _06418_ _06419_ _06420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_139_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11635_ _01068_ _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_53_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11578__A1 _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17142_ _00212_ clknet_leaf_128_clk channels.atk_dec2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_24_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14354_ _06219_ _06227_ _06352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11566_ _03639_ _03680_ _03683_ _00414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_80_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13305_ _05309_ _05310_ _05311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__10250__A1 _01508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17073_ _00143_ clknet_leaf_119_clk net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10517_ _02504_ _02777_ _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14285_ _03345_ _05853_ _06284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11497_ channels.freq1\[4\] _03633_ _03634_ _03635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16024_ _07822_ _07827_ _07904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13236_ _05067_ _05071_ _05242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_110_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10448_ _02685_ _02628_ _02703_ _02708_ _02709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_13167_ _05067_ _05071_ _05172_ _05173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10379_ _02629_ _02631_ _02639_ _02640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_23_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12118_ channels.accum\[3\]\[7\] _04141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13098_ _03270_ _04240_ _04816_ _05104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_88_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16926_ tt_um_rejunity_sn76489.control_noise\[0\]\[0\] _00993_ _00877_ _00994_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12049_ _04100_ _00480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11502__A1 _02326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16857_ _02707_ _03742_ _03128_ _02847_ _00945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_46_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15808_ _06858_ _07690_ _07704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16788_ _00895_ _00897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13255__A1 _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09550__I _01904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15739_ _07653_ _07654_ _00616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13072__I _05077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09260_ channels.lfsr\[3\]\[15\] _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09191_ channels.lfsr\[2\]\[7\] _01633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_90_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17409_ _00479_ clknet_leaf_158_clk channels.adsr_state\[3\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_173_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11569__A1 channels.freq3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14507__A1 _06298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08737__A2 _01105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09725__I channels.pw1\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08975_ _01437_ _01438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__16680__A1 _08419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14787__B _06775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09162__A2 _01592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16558__I _01752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15235__A2 _07149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13246__A1 _05069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09527_ _01762_ _01844_ _01848_ channels.pw2\[1\] _01916_ _01917_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_79_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14994__A1 filters.filt_3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09458_ _01000_ _01839_ _01849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_13_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13549__A2 _05454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14746__A1 _06403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09389_ _01786_ _01787_ _01788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_49_Left_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11420_ _03578_ _01571_ _03588_ _00363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_173_3593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11351_ _01585_ _03534_ _03544_ _03545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_22_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_134_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10302_ _02555_ _02562_ _02563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14070_ _06065_ _06069_ _06071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11282_ _02316_ _03484_ _03488_ _00325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_104_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16242__B _07700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09925__A1 channels.sus_rel2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13021_ _05025_ _05007_ _05026_ _05027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_10233_ _02423_ _02474_ _02489_ _02493_ _02494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__10535__A2 _02754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10164_ _01097_ _01098_ channels.pw2\[7\] _02425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XPHY_EDGE_ROW_58_Left_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_17760_ _00830_ clknet_leaf_70_clk tt_um_rejunity_sn76489.latch_control_reg\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14972_ _06942_ _06943_ _06944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10095_ _02358_ _02359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10299__A1 _01328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_6_clk_I clknet_5_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16711_ _03710_ _08446_ _08448_ _00794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13923_ _04483_ _04818_ _05925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17691_ _00761_ clknet_leaf_216_clk channels.lfsr\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_210_clk clknet_5_20__leaf_clk clknet_leaf_210_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__15226__A2 _07187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16642_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[3\] tt_um_rejunity_sn76489.tone\[0\].gen.counter\[2\]
+ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[1\] tt_um_rejunity_sn76489.tone\[0\].gen.counter\[0\]
+ _08391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__08900__A2 _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13854_ _05752_ _05755_ _05857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_69_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12805_ _04799_ _04810_ _04811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_69_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16573_ _08314_ _08351_ _00753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14985__A1 filters.high\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13785_ _05696_ _05786_ _05788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11405__I _01089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10997_ _03221_ _03222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_44_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15524_ _03264_ _07463_ _07464_ _03218_ _07465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_26_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12736_ _04198_ _04742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_127_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12460__A2 _04327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_67_Left_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_128_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15455_ _07398_ _07400_ _07401_ _07402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_12667_ _04663_ _04670_ _04671_ _04672_ _04673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__14716__I _06067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13620__I _05145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14406_ _05543_ _06403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11618_ _03664_ _03712_ _03717_ _00432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_53_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15386_ _07328_ _07337_ _07338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12598_ _04598_ _04602_ _04603_ _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_108_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17125_ _00195_ clknet_leaf_117_clk channels.pw2\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14337_ _06211_ _06212_ _06335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11549_ _03651_ _03671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10774__A2 _02840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17056_ _00126_ clknet_leaf_89_clk filters.filt_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14268_ _06265_ _06266_ _06267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_40_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16007_ _07853_ _07886_ _07887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_59_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13219_ _05224_ _05217_ _05225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_59_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14199_ _06114_ _06198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_57_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09545__I _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08760_ _01239_ _00048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_178_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16909_ channels.exp_counter\[3\]\[3\] _00984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__16378__I _08194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08691_ _01152_ _01175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_135_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15217__A2 _02029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_201_clk clknet_5_23__leaf_clk clknet_leaf_201_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_178_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13243__A4 _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09312_ _01632_ _01729_ _01731_ _01636_ _00108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_24_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12451__A2 _04390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14991__A4 channels.sample2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09243_ channels.lfsr\[3\]\[13\] _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15231__B _07086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14728__A1 _06720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09174_ channels.lfsr\[3\]\[3\] _01619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11411__B1 _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_151_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput27 net27 bus_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_112_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10517__A2 _02777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15456__A2 _06983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08958_ _01321_ _01422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__15406__B _07356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08889_ _01349_ _01358_ _01359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10920_ channels.sample2\[10\] _03156_ _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_169_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_158_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10851_ _03085_ _03103_ _03104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_66_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_175_3633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13570_ _05569_ _05574_ _05575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_66_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12442__A2 _04447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10782_ _03027_ _03036_ _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_137_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12521_ _04523_ _04524_ _04526_ _04527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__14719__A1 _06689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_137_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13440__I _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15240_ _07197_ _07201_ _07202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12452_ _03254_ _04225_ _04376_ _04458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_11403_ _03578_ _01515_ _03579_ _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15171_ _07112_ _07136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_90_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13942__A2 _05943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12383_ _03286_ _04195_ _04389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_133_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14122_ _06107_ _06121_ _06122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11334_ _03515_ _03522_ _03528_ _00337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_160_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16341__B1 _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14053_ _06045_ _06053_ _06054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_162_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11265_ _03474_ _03475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11828__C _01170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11705__A1 channels.sus_rel3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11705__B2 channels.sus_rel2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13004_ _04462_ _05006_ _05007_ _05010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_24_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10216_ _02438_ _02442_ _02477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_37_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11196_ filters.high\[11\] _03410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_37_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10147_ channels.pw1\[9\] _01251_ _02408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11469__B1 _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17743_ _00813_ clknet_leaf_54_clk tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14955_ _06911_ _06912_ _06927_ _06928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10078_ filters.cutoff_lut\[16\] _02341_ _02342_ _02346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_168_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13906_ _05820_ _05906_ _05907_ _05908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_17674_ _00744_ clknet_leaf_81_clk tt_um_rejunity_sn76489.tone\[2\].gen.counter\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14886_ _06768_ _06853_ _06865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_43_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13837_ _05834_ _05839_ _05840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_16625_ _01663_ _08384_ _08385_ _01665_ _00771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08980__S1 _01164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16556_ _08323_ _08335_ _08334_ _08337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_128_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13768_ _05683_ _05702_ _05771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_70_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10444__A1 _01162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15507_ _03194_ _04189_ _07446_ _07449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_12719_ _04458_ _04459_ _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_45_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16487_ _08274_ _08277_ _08278_ _08279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xclkbuf_0_clk clk clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13699_ _05683_ _05702_ _05703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_26_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15438_ _07383_ _07384_ _07385_ _07386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_26_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15369_ filters.high\[20\] _07310_ _07223_ _07323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_96_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09062__A1 _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17108_ _00178_ clknet_leaf_111_clk channels.sus_rel1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09930_ _01818_ _02242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17039_ _00109_ clknet_leaf_223_clk channels.lfsr\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09861_ channels.ctrl_reg2\[0\] _02195_ _02189_ _02196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_111_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08812_ _01284_ _01285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_212_clk_I clknet_5_20__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09792_ _02110_ _02142_ _02145_ _00178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13449__A1 _05444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08743_ channels.exp_counter\[1\]\[1\] _01105_ _01225_ _01220_ _01226_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_139_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08674_ _01157_ _01158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12672__A2 _04675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_227_clk_I clknet_5_17__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_152_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10089__C _02354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_5_4__f_clk_I clknet_3_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_153_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09226_ _01658_ _01659_ _01663_ _01651_ _00090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_91_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_170_3530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_170_3541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09157_ _01201_ _01604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_146_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_131_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09088_ _01541_ _01542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_169_Right_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__17319__D _00389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11050_ _03272_ _03273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10001_ _02290_ _02292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_129_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_129_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14740_ _06703_ _06731_ _06732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_11952_ channels.env_counter\[2\]\[4\] _04030_ _04031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_28_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10123__B1 _01286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08867__A1 _01327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16929__A2 _00993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13860__A1 _05547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10903_ _03147_ _02932_ _03148_ _00286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14671_ _06580_ _06588_ _06666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11883_ _03961_ _03969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16410_ _08217_ _08218_ _08211_ _00723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13622_ _05231_ _05624_ _05626_ _04473_ _05627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_17390_ _00460_ clknet_leaf_148_clk channels.env_counter\[2\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10834_ _03028_ _02939_ _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13612__A1 _05484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12415__A2 _04420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16341_ _01218_ _01255_ _01258_ channels.exp_counter\[0\]\[0\] _08171_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_13553_ _05459_ _05525_ _05558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08714__S1 _01172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10765_ _02987_ _03006_ _03020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12504_ _04396_ _04510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16272_ filters.sample_buff\[12\] _07742_ _08130_ spi_dac_i.spi_dat_buff_0\[8\] spi_dac_i.spi_dat_buff_0\[9\]
+ _08127_ _08133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_109_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13484_ _05484_ _05489_ _05490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_70_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10696_ _02602_ _02623_ _02953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15223_ _07183_ _07184_ _07185_ _07186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_12435_ filters.filter_step\[2\] _03181_ filters.filter_step\[0\] _04441_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_0_65_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09044__A1 _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_164_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09595__A2 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15154_ _06913_ _07119_ _07120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_39_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12366_ _04371_ _04372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_106_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_136_Right_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15097__I _06913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14105_ _06042_ _06054_ _06104_ _06105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_11317_ _02333_ _03516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15085_ net31 _05043_ _05048_ _07053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__13679__A1 _05591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12297_ _04301_ _04302_ _04303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_91_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14036_ _04801_ _04923_ _06037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_91_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11248_ filters.high\[14\] _03235_ _03459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_129_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12351__A1 _04252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11179_ filters.low\[10\] _03394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16093__A2 _07942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15987_ spi_dac_i.counter\[0\] _07725_ _07868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13345__I _05350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17726_ _00796_ clknet_leaf_60_clk tt_um_rejunity_sn76489.control_tone_freq\[2\]\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_145_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14938_ _04558_ _04690_ _06912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08858__A1 _01327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_17657_ _00727_ clknet_leaf_52_clk tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14869_ filters.band\[25\] _06820_ _06811_ _06850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15560__I _01932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16608_ _01580_ _08376_ _08379_ _01595_ _00760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_9_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17588_ _00658_ clknet_leaf_44_clk spi_dac_i.spi_dat_buff_1\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_147_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16539_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[9\] tt_um_rejunity_sn76489.tone\[1\].gen.counter\[8\]
+ _08320_ _08321_ _08322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_45_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_93_clk_I clknet_5_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09011_ _01471_ _01472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10209__I channels.pw2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_103_Right_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09913_ _02185_ _02227_ _02230_ _00214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_151_clk_I clknet_5_29__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09844_ channels.pw2\[8\] _02182_ _02176_ _02183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_176_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_146_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09775_ _02124_ _02134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_13_Left_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_166_clk_I clknet_5_25__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08726_ _01179_ _01208_ _01209_ _01188_ _01210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_69_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08657_ _01140_ _01141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_96_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_46_clk_I clknet_5_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08588_ _01103_ _01104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_113_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14086__I _05990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13070__A2 _05075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10550_ _02522_ _02622_ _02810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09209_ channels.lfsr\[3\]\[8\] _01649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_88_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_104_clk_I clknet_5_13__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10481_ _02627_ _02640_ _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_161_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09908__I _02226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12220_ _04225_ _04226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_121_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10187__A3 channels.pw2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08785__B1 _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12151_ _04157_ _00525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11102_ _03305_ _03322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_119_clk_I clknet_5_26__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12082_ channels.env_counter\[0\]\[9\] _04120_ _04122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14322__A2 _06027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15910_ _07791_ _07792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_11033_ filters.low\[1\] _03187_ _03256_ _03206_ _03257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_159_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16890_ _01583_ _03739_ _00973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_21_1168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_1225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15841_ spi_dac_i.counter\[0\] _07726_ _07727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10895__A1 channels.sample2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15822__A2 _07640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12984_ _04987_ net52 _04990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_15772_ _06758_ _07677_ _07678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_99_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17511_ _00581_ clknet_leaf_27_clk filters.high\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11935_ _04009_ _04015_ _04016_ _04017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__08935__S1 _01163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14723_ _06703_ _06716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15380__I _07332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17442_ _00512_ clknet_leaf_147_clk channels.accum\[3\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14654_ _06640_ _06642_ _06648_ _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_135_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11866_ channels.env_vol\[0\]\[2\] _03942_ _03955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13605_ _05478_ _05608_ _05609_ _05610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10817_ _03063_ _03070_ _03071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_14585_ _06421_ _06422_ _06581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_17373_ _00443_ clknet_leaf_210_clk channels.env_vol\[0\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11797_ _03887_ _03888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13061__A2 _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16324_ _03743_ _08158_ _08161_ _00694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_83_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13536_ filters.band\[0\] _05540_ _05541_ _05542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10748_ _03000_ _03003_ _03004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_165_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16255_ _08116_ _08122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10029__I _02293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13467_ _05470_ _05471_ _05472_ _05473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_10679_ _02885_ _02934_ _02935_ _02936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_129_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15206_ _07146_ _07149_ _07169_ _07170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09568__A2 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12418_ _04292_ _04208_ _04424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16186_ _07995_ _08060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13398_ _05403_ _05379_ _05404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_112_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15137_ _07074_ _07075_ _07103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12349_ _04325_ _04355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_50_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08871__S0 _01145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_71_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15068_ _07001_ _07003_ _07027_ _07006_ _07036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__15510__A1 _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14019_ _06011_ _06019_ _06020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_156_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16066__A2 _07914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10886__A1 channels.sample3\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09560_ channels.atk_dec1\[2\] _01948_ _01949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_175_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08511_ _01028_ _01038_ _01039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_19_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17709_ _00779_ clknet_leaf_228_clk channels.lfsr\[0\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_69_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09491_ _01881_ _01882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_19_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_136_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15577__A1 _01927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_102_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15329__A1 _07277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09728__I _01062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_rebuffer28_I _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09103__S1 _01480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12154__I _04159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16070__B _07721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_21_Left_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_109_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09827_ _02162_ _02170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_126_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14068__A1 _03314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15804__A2 _07640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09758_ channels.ctrl_reg1\[7\] _02117_ _02120_ _02122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_154_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08709_ channels.exp_periods\[2\]\[4\] _01193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09689_ _02060_ _02071_ _02072_ _00148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_167_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11720_ channels.atk_dec3\[6\] _01439_ _03783_ channels.atk_dec2\[6\] _01291_ channels.atk_dec1\[6\]
+ _03811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_68_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output19_I net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11651_ _02839_ _03742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_30_Left_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14240__A1 filters.band\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10602_ _02536_ _02622_ _02861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14370_ _06358_ _06367_ _06368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_181_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11582_ _03675_ _03687_ _03693_ _00420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_135_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13321_ _04395_ _04375_ _05327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10533_ _02744_ _02762_ _02793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08470__A2 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16040_ _07873_ _07919_ _07920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13252_ _04199_ _04862_ _05258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_150_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10464_ _02717_ _02718_ _02725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12203_ _04206_ _04208_ _04209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12554__A1 _04528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11357__A2 _03549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13183_ _05182_ _05184_ _05188_ _05189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_10395_ _02655_ _02644_ _02630_ _02656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_103_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12134_ channels.accum\[3\]\[15\] _04149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12065_ _04021_ _04105_ _04111_ _00485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16942_ _00021_ clknet_leaf_221_clk channels.lfsr\[3\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11016_ _01069_ _03227_ _03240_ _03241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_159_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16873_ _03746_ _00959_ _00960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_159_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15824_ _04189_ _04158_ _07713_ _00642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xclkbuf_5_24__f_clk clknet_3_6_0_clk clknet_5_24__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_99_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12967_ _04964_ _04961_ _04973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_35_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15755_ _07665_ _07666_ _00620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11918_ _03834_ _03987_ _04000_ _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_14706_ _06688_ _06700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_169_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15686_ _07608_ _07614_ _07573_ _00603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_12898_ _04902_ _04903_ _04904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_47_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17425_ _00495_ clknet_leaf_130_clk channels.env_counter\[0\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_157_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14637_ _06585_ _06586_ _06632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_51_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11849_ _01087_ _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__14231__A1 _06197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14568_ _04355_ _05775_ _06442_ _06564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_17356_ _00426_ clknet_leaf_172_clk channels.pw3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12793__A1 _04787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16307_ channels.env_counter\[3\]\[9\] _08151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10982__I _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13519_ _05494_ _05524_ _05525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_67_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14499_ _06495_ _06496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_17287_ _00357_ clknet_leaf_190_clk channels.accum\[2\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_141_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16238_ spi_dac_i.spi_dat_buff_1\[10\] _07870_ _08098_ _08110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_125_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15731__A1 _05969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16169_ _08042_ _08043_ _08044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09410__A1 _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09961__A2 _01842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08991_ _01451_ _01452_ _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_142_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14298__B2 _06285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_143_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09612_ _01881_ _01999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_3_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09543_ _01931_ _01932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09021__S0 _01138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09474_ _01748_ _01844_ _01848_ channels.pw2\[0\] _01864_ _01865_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_149_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_119_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16278__A2 _07742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10180_ _02428_ channels.pw2\[4\] _01097_ _02441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__12839__A2 _04796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_180_3724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13870_ _05747_ _05657_ _05849_ _05872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_9_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09921__I _02226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12821_ _04822_ _04823_ _04826_ _04827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_119_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13264__A2 _05268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15540_ _07472_ _07473_ _07479_ _07480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_12752_ _04713_ _04758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_178_3686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11703_ _03533_ _03787_ _03790_ _03793_ _03794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_15471_ filters.low\[29\] _07416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_12683_ _04685_ _04687_ _04689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_167_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14422_ _06322_ _06323_ _06419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_17210_ _00280_ clknet_leaf_93_clk channels.sample3\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11634_ _03727_ _03728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_182_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17141_ _00211_ clknet_leaf_127_clk channels.atk_dec2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_154_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14353_ _06221_ _06226_ _06351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_181_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11565_ channels.freq3\[0\] _03681_ _03682_ _03683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_42_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09640__A1 channels.sus_rel2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13304_ _03285_ _04194_ _05106_ _05310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_17072_ _00142_ clknet_leaf_113_clk net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10516_ _02776_ _02777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_134_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14284_ _06278_ _06282_ _06283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__10250__A2 _02381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11496_ _03516_ _03634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16023_ _07899_ _07902_ _07903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_150_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13235_ _05207_ _05225_ _05240_ _05241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_10447_ _02704_ _02707_ _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_110_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13166_ _05068_ _05070_ _05172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_10378_ _02509_ _02569_ _02638_ _02639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_62_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12117_ _04140_ _00508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13097_ _04883_ _04885_ _05103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_88_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16925_ _03490_ _00922_ _03519_ _00993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_12048_ channels.adsr_state\[3\]\[1\] _04100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_88_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16856_ _03746_ _00941_ _00943_ _00944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_49_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15807_ _07702_ _07703_ _00635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09459__A1 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16787_ _00895_ _00896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_149_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13255__A2 _05260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13999_ _05998_ _05958_ _05999_ _06000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_66_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15738_ _03329_ _07643_ _07644_ _07654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_141_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15669_ filters.sample_buff\[11\] _07592_ _07599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17408_ _00478_ clknet_leaf_129_clk channels.env_counter\[1\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09190_ _01628_ _01611_ _01632_ _01627_ _00085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_172_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17339_ _00409_ clknet_leaf_103_clk channels.freq2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12518__A1 _03273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08974_ _01427_ _01428_ _01437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_89_Right_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09698__A1 channels.freq1\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11048__I _03270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13246__A2 _04750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14443__A1 _04453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09526_ _01913_ _01914_ _01915_ _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_149_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14994__A2 channels.sample3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09457_ _01847_ _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_8_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_98_Right_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_164_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09388_ net1 _01787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_53_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_3594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11350_ _02847_ _03543_ _03544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_22_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10301_ _02561_ _02562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_132_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11281_ filters.cutoff_lut\[8\] _03483_ _03485_ _03488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_131_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13182__A1 _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13020_ _04996_ _04998_ _05000_ _05026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_131_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10232_ _02459_ _02490_ _02492_ _02493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__17057__D _00127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10163_ _02423_ _02424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_5_Left_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__16749__I _00867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14971_ _01768_ channels.sample3\[1\] _06943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10094_ _02357_ _02358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14682__A1 _04453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16710_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[4\] _08447_ _08318_ _08448_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13922_ _04396_ _05731_ _05924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17690_ _00760_ clknet_leaf_213_clk channels.lfsr\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16641_ _01720_ _08375_ _08378_ _08390_ _00782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_18_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13853_ _05852_ _05855_ _05856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_57_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12804_ _04808_ _04809_ _04810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16572_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[4\] _08347_ _08349_ _08350_
+ _08351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_13784_ _05696_ _05786_ _05787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14985__A2 _06955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10996_ _03220_ _03221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_96_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15523_ channels.sample3\[1\] _07452_ _07464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12735_ _04184_ _04740_ _04741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_1307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09861__A1 channels.ctrl_reg2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12460__A3 _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15454_ _07398_ _07400_ _07240_ _07401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_61_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12666_ _04657_ _04659_ _04672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12748__A1 _04286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11617_ channels.pw2\[2\] _03713_ _03714_ _03717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14405_ _03361_ _06080_ _06402_ _06187_ _00534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_182_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09613__A1 channels.freq3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12597_ _04353_ _04297_ _04599_ _04601_ _04603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_15385_ _07327_ _06836_ _07337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_108_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09613__B2 channels.ctrl_reg3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17124_ _00194_ clknet_leaf_118_clk channels.pw2\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_41_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11420__A1 _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11548_ _03657_ _03670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14336_ _06223_ _06224_ _06333_ _06334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_80_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17055_ _00125_ clknet_leaf_90_clk filters.filt_1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14267_ _05440_ _06096_ _06266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11479_ _00131_ _01033_ _01029_ _03623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_151_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16006_ _07791_ _07799_ _07886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13218_ _05222_ _05223_ _05224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_59_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14198_ _06195_ _06196_ _06197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_59_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12252__I _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13149_ _05111_ _05112_ _05155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__11296__C _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14673__A1 _04806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11487__A1 _02308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16908_ _00983_ _00849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_174_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08690_ _01173_ _01174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_139_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16839_ tt_um_rejunity_sn76489.clk_counter\[1\] _00928_ _03729_ _00931_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_75_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09311_ _01625_ _01729_ _01731_ _01630_ _00107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09242_ channels.lfsr\[1\]\[13\] _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_173_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10462__A2 _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14728__A2 _06712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12739__A1 _04732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09173_ channels.lfsr\[1\]\[3\] _01618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09080__A2 _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer10_I _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09736__I _02106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13164__A1 _05121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput28 net28 bus_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_141_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12911__A1 _04853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16653__A2 _08267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08957_ _01408_ _01409_ _01420_ _01421_ _00063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_76_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11707__S _03784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11478__A1 _03612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08888_ _01351_ _01357_ _01358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09540__B1 net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11506__I _01779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_158_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10850_ _03086_ _03102_ _03103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_175_3623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09509_ _01856_ _01846_ _01900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_52_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_175_3634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10781_ _03029_ _03035_ _03036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_177_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12520_ _03317_ _04525_ _04164_ _04526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_93_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11650__A1 _01933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14719__A2 _06712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_117_Right_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_136_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12451_ _04366_ _04390_ _04457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_81_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_164_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11402_ channels.accum\[2\]\[15\] _03571_ _03579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10205__A2 channels.pw2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15170_ net56 _07122_ _07134_ _07135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_133_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12382_ _04253_ _04388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_62_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14121_ _06115_ _06120_ _06121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11333_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[3\] _03523_ _03517_ _03528_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_10_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_21__f_clk_I clknet_3_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14052_ _06048_ _06052_ _06053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_104_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11264_ _03473_ _03474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_31_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12902__A1 _04852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13003_ _04996_ _05001_ _05009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10215_ _01541_ _02433_ _02452_ _01533_ _02476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_11195_ filters.sample_filtered\[11\] _03409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_24_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_37_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10146_ _02390_ channels.pw2\[9\] _02397_ _02407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_17742_ _00812_ clknet_leaf_54_clk tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12800__I _04805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10077_ _02326_ _02340_ _02345_ _00263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14954_ _06926_ _06927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09381__I _01779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13905_ _05821_ _05822_ _05907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_17673_ _00743_ clknet_leaf_59_clk tt_um_rejunity_sn76489.tone\[2\].gen.counter\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14885_ _06862_ _06863_ _06864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_195_clk clknet_5_23__leaf_clk clknet_leaf_195_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16624_ _01657_ _08384_ _08385_ _01660_ _00770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_134_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13836_ _05835_ _05838_ _05839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_173_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_175_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16555_ _08323_ _08334_ _08335_ _08336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_174_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15332__B _06899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_174_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13767_ _05686_ _05701_ _05770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10979_ _03203_ _03204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_168_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_174_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15506_ _07447_ _07448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_85_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12718_ _04458_ _04459_ _04724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16486_ _08261_ _08276_ _08275_ _08278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_57_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13698_ _05686_ _05701_ _05702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_85_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15437_ _07372_ _06765_ _07385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12247__I _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12649_ _04653_ _04654_ _04598_ _04655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__15383__A2 _06919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15368_ _07315_ _07321_ _07322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_142_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_96_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09062__A2 _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17107_ _00177_ clknet_leaf_112_clk channels.sus_rel1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14319_ _06205_ _06206_ _06317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15299_ filters.high\[14\] _06955_ _07258_ _07259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13146__A1 _05142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_141_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17038_ _00108_ clknet_leaf_223_clk channels.lfsr\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_74_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09860_ _02193_ _02195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08811_ _01248_ channels.clk_div\[1\] _01284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09791_ channels.sus_rel1\[1\] _02143_ _02138_ _02145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15507__B _07446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13449__A2 _05454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14646__A1 _04576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08742_ _01217_ _01224_ _01225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__14110__A3 _05106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09522__B1 _01842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08673_ _01156_ _01157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10132__A1 channels.pw1\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_186_clk clknet_5_22__leaf_clk clknet_leaf_186_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_17_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09825__A1 channels.freq2\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13541__I _05543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11632__A1 _03677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09225_ _01660_ _01661_ _01652_ _01662_ _01643_ _01644_ _01663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_174_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_170_3531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_170_3542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09156_ channels.lfsr\[3\]\[1\] _01603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_32_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_5_clk_I clknet_5_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09053__A2 _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11396__B1 _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_86_Left_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_131_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09087_ channels.accum\[0\]\[19\] channels.accum\[1\]\[19\] channels.accum\[2\]\[19\]
+ channels.accum\[3\]\[19\] _01495_ _01496_ _01541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_102_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_110_clk clknet_5_15__leaf_clk clknet_leaf_110_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_131_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_168_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10000_ _02290_ _02291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09989_ _02254_ _02284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_157_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_129_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_5_5__f_clk clknet_3_1_0_clk clknet_5_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_129_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_95_Left_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11951_ _04011_ _04030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10123__A1 channels.ctrl_reg2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_177_clk clknet_5_18__leaf_clk clknet_leaf_177_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10123__B2 channels.ctrl_reg1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10902_ channels.sample2\[3\] _03143_ _03148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_168_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14670_ _06580_ _06588_ _06665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11882_ _02752_ _03538_ _03967_ _03968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_98_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13621_ _05625_ _05626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10833_ _03074_ _03076_ _03086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_79_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13612__A2 _05489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16340_ _03981_ _08165_ _08170_ _00701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08545__I net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13552_ _05494_ _05524_ _05557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10764_ _02990_ _03005_ _03019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12503_ _04398_ _04507_ _04508_ _04509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_109_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16271_ _08129_ _08132_ _00670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13483_ _05485_ _05486_ _05488_ _05489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_10695_ _02901_ _02902_ _02904_ _02952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_124_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_164_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12434_ _04381_ _04439_ _04440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_15222_ _01748_ channels.sample1\[10\] _07185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_168_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11387__B1 _01420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12365_ _04314_ _04371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15153_ _07095_ _07118_ _07119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_106_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_101_clk clknet_5_13__leaf_clk clknet_leaf_101_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_26_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_39_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11316_ _02298_ _03515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_14104_ _06026_ _06041_ _06104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_10_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16865__A2 _02455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15084_ filters.low\[6\] _07051_ _07052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_121_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12296_ _04207_ _04302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14035_ _06030_ _06035_ _06036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_91_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10315__I _02575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11247_ _03455_ _03226_ _03457_ _03458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_38_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11178_ _03242_ _03393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_52_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14628__A1 _05909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10129_ _01272_ _02390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15986_ _07729_ _07867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_175_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17725_ _00795_ clknet_leaf_59_clk tt_um_rejunity_sn76489.control_tone_freq\[2\]\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_136_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10114__A1 channels.ctrl_reg1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14937_ filters.low\[0\] _06911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_168_clk clknet_5_25__leaf_clk clknet_leaf_168_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11146__I _03362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17656_ _00726_ clknet_leaf_52_clk tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14868_ _06804_ _06848_ _06849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_58_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16607_ _08378_ _08379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13819_ _04893_ _05518_ _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15062__B _07030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09807__A1 _02155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17587_ _00657_ clknet_leaf_45_clk spi_dac_i.spi_dat_buff_1\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13361__I _05187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14799_ _06784_ _06786_ _00544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_161_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16538_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[7\] tt_um_rejunity_sn76489.tone\[1\].gen.counter\[6\]
+ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[5\] tt_um_rejunity_sn76489.tone\[1\].gen.counter\[4\]
+ _08321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__11614__A1 _03710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16469_ _08237_ _08263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09010_ _01468_ _01470_ _01471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_54_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_83_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_76_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15108__A2 channels.sample1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09912_ channels.sus_rel2\[1\] _02228_ _02224_ _02230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09843_ _02180_ _02182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_146_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09774_ _02124_ _02133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_146_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08725_ _01187_ channels.exp_periods\[3\]\[1\] _01209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10105__A1 _02366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_159_clk clknet_5_28__leaf_clk clknet_leaf_159_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__15751__I _07635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08656_ _01139_ _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_178_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16241__B1 _08111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_124_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_138_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08587_ _01102_ _01100_ _01103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__16792__A1 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11605__A1 _03675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16919__I0 _00966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09208_ channels.lfsr\[1\]\[8\] _01648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10480_ _02626_ _02739_ _02740_ _02741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_63_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09139_ _01581_ _01587_ _01588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__08785__A1 _01086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12150_ channels.accum\[3\]\[23\] _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08785__B2 channels.ring_outs\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11101_ filters.sample_filtered\[5\] _03320_ _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12081_ _04047_ _04119_ _04121_ _00491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_124_1164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09924__I _02154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11032_ _03255_ _03256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_34_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15840_ _07725_ _07726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_95_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15771_ _07663_ _07677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12983_ _04987_ _04988_ _04989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_17510_ _00580_ clknet_leaf_27_clk filters.high\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14722_ _04161_ _06714_ _06715_ _00538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_99_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11934_ _03880_ _03874_ _04016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__15035__A1 _06983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17441_ _00511_ clknet_leaf_163_clk channels.accum\[3\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14653_ _06643_ _06646_ _06647_ _06648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_157_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11865_ _03747_ _03953_ _03954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_68_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13604_ _05479_ _05480_ _05609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_17372_ _00442_ clknet_leaf_208_clk channels.env_vol\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10816_ _03064_ _03069_ _03070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_55_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11796_ channels.env_counter\[0\]\[3\] channels.env_counter\[1\]\[3\] channels.env_counter\[2\]\[3\]
+ channels.env_counter\[3\]\[3\] _03886_ _01166_ _03887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_14584_ _06577_ _06578_ _06579_ _06580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_6_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16323_ channels.env_vol\[1\]\[0\] _08160_ _08161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_166_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13535_ _03721_ _05541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_131_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10747_ _03001_ _03002_ _03003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_83_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_211_clk_I clknet_5_20__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16254_ _07597_ _08121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13466_ _04317_ _04752_ _05472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10678_ _02888_ _02930_ _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15205_ _07164_ _07168_ _07169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_93_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12417_ _04340_ _04345_ _04422_ _04423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16185_ _07811_ _07904_ _07911_ _08059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_51_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13397_ _05391_ _05401_ _05402_ _05403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_65_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__16838__A2 _03731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15136_ _07073_ _07102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12348_ _04353_ _04354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_121_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_226_clk_I clknet_5_20__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08871__S1 _01159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12279_ _04249_ _04284_ _04285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_71_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15067_ _07030_ _07035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_120_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15510__A2 _03204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09834__I _02174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14018_ _06014_ _06018_ _06019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__12260__I _04265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15969_ _07801_ _07791_ _07850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08510_ _00132_ _01035_ _01037_ _01038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_17708_ _00778_ clknet_leaf_229_clk channels.lfsr\[0\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09490_ _01850_ _01840_ _01881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_72_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15504__C _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08700__A1 _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17639_ _00709_ clknet_leaf_208_clk channels.ch3_env\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__14187__I _06186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16774__A1 _03499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13588__A1 _04848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_102_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09256__A2 _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10810__A2 _02872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_148_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_165_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10326__A1 _01598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09826_ _02131_ _02163_ _02169_ _00188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_126_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14068__A2 _06067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09757_ _01814_ _02116_ _02121_ _00167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13815__A2 _05723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08708_ channels.exp_periods\[0\]\[4\] channels.exp_periods\[1\]\[4\] _01178_ _01192_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_154_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_169_Left_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09688_ net29 _01909_ _02036_ _02072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15017__A1 filters.filt_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08639_ _01130_ _00036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__16765__A1 _01806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11650_ _01933_ _03741_ _00440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09247__A2 _01659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10601_ _02594_ _02500_ _02860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11581_ channels.freq3\[6\] _03688_ _03690_ _03693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09919__I _02149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13320_ _04323_ _04489_ _05326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10532_ _02767_ _02778_ _02791_ _02792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12003__A1 _03925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10463_ _02654_ _02716_ _02724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13251_ _04266_ _05256_ _05257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_178_Left_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_122_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12202_ _04207_ _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13182_ _04401_ _05187_ _05188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_10394_ _02598_ _02655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10565__A1 _02607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12133_ _04148_ _00516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_130_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12064_ channels.env_counter\[0\]\[2\] _04108_ _04111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16941_ _00020_ clknet_leaf_221_clk channels.lfsr\[3\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11015_ filters.hp _03236_ _03237_ filters.bp _03239_ _03240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_16872_ _00941_ _00950_ _00959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_102_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15256__A1 _03422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08930__A1 _01389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15823_ _03735_ _07628_ _07713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_5_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11817__A1 _03905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15754_ _03394_ _07656_ _07657_ _07666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_133_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12966_ _04965_ _04970_ _04971_ _04972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_87_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14705_ _06602_ _06699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_11917_ _03989_ _03990_ _03999_ _04000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_15685_ _07450_ _07612_ _07613_ _07614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12897_ _03316_ _04163_ _04450_ _04903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_47_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17424_ _00494_ clknet_leaf_148_clk channels.env_counter\[0\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14636_ _06585_ _06586_ _06631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_47_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11848_ _03938_ _03939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_172_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_150_clk_I clknet_5_29__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14231__A2 _06229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_64_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17355_ _00425_ clknet_leaf_95_clk channels.pw3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12242__A1 _04233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14567_ _06561_ _06562_ _06563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11779_ _03804_ _03869_ _03870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16306_ _08150_ _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08997__A1 _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13518_ _05497_ _05523_ _05524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13990__A1 _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_30_clk_I clknet_5_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17286_ _00356_ clknet_leaf_158_clk channels.accum\[2\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14498_ _06390_ _06394_ _06495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_3_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16237_ spi_dac_i.spi_dat_buff_1\[9\] _07834_ _08096_ _08108_ _08109_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_42_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13449_ _05444_ _05454_ _05455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_2_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_165_clk_I clknet_5_25__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16168_ _08041_ _08038_ _08039_ _08043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_23_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_45_clk_I clknet_5_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15119_ _07029_ _07086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_103_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08990_ channels.freq2\[11\] _01279_ _01292_ channels.freq1\[11\] _01452_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_16099_ _07969_ _07972_ _07976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14298__A2 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_143_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_143_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09611_ channels.pw2\[4\] _01996_ _01997_ channels.freq2\[12\] _01998_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08921__B2 channels.freq1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_160_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_103_clk_I clknet_5_13__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09542_ _01087_ _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_167_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09021__S1 _01480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16747__A1 _01806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09473_ _01852_ _01858_ _01863_ _01864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_116_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_84_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_90_clk clknet_5_12__leaf_clk clknet_leaf_90_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_149_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_118_clk_I clknet_5_26__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12233__A1 _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08988__A1 _01442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12536__A2 _04541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17608__D _00678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_30__f_clk clknet_3_7_0_clk clknet_5_30__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_30_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_160_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14289__A2 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11509__I _03641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_180_3725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09809_ _02137_ _02158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_92_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12820_ _03254_ _04225_ _04825_ _04826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_119_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12751_ _04738_ _04755_ _04756_ _04757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_81_clk clknet_5_9__leaf_clk clknet_leaf_81_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_178_3687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11702_ _03791_ _03792_ _03793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15470_ filters.low\[28\] _06766_ _07415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_38_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12682_ _04687_ _04685_ _04688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_155_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14213__A2 _05075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14421_ _06320_ _06321_ _06418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11633_ _01092_ _01093_ _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_181_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_139_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17140_ _00210_ clknet_leaf_128_clk channels.atk_dec2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_92_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14352_ _06348_ _06349_ _06350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11564_ _03651_ _03682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13303_ _03300_ _04276_ _04879_ _05309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_17071_ _00141_ clknet_leaf_119_clk net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10515_ _02775_ _02776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11495_ _03624_ _03633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14283_ _06279_ _06175_ _06281_ _06282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_134_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15713__A2 _07632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16022_ _07900_ _07901_ _07902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__13724__A1 _05630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12527__A2 _04528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13234_ _05228_ _05234_ _05239_ _05240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_10446_ _02706_ _02707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13165_ _05117_ _05169_ _05170_ _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_10377_ _02637_ _02638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_62_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12116_ channels.accum\[3\]\[6\] _04140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13096_ _04886_ _04890_ _05102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_137_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16924_ _00992_ _00856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12047_ _04099_ _00479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_88_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08903__A1 _01337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16855_ _03536_ _03128_ _03131_ _00942_ _00943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_88_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15806_ _07373_ _07694_ _07695_ _07703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_49_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16786_ _00879_ _00894_ _00895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13998_ _05905_ _05935_ _05999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_66_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15737_ _06184_ _07652_ _07653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_87_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12949_ _04475_ _04482_ _04955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_133_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_72_clk clknet_5_14__leaf_clk clknet_leaf_72_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_153_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15668_ _07597_ _07598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_34_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17407_ _00477_ clknet_leaf_130_clk channels.env_counter\[1\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14619_ _06356_ _06614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_157_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16881__S _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15599_ filters.sample_buff\[6\] _07461_ _07523_ _07534_ _07535_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_29_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17338_ _00408_ clknet_leaf_103_clk channels.freq2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09631__A2 net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17269_ _00339_ clknet_leaf_153_clk channels.adsr_state\[0\]\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_178_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08973_ _01298_ _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_162_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09525_ channels.sus_rel3\[1\] _01859_ _01861_ channels.pw2\[9\] _01915_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_149_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_63_clk clknet_5_11__leaf_clk clknet_leaf_63_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_66_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09456_ _01826_ _01846_ _01847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_149_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09387_ net2 _01786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_19_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_173_3595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10300_ _01328_ _02558_ _02560_ _02561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_134_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11280_ _02314_ _03484_ _03487_ _00324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_134_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09386__A1 net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10231_ _02460_ _02491_ _01469_ _02492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13182__A2 _05187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12623__I _04420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11812__S0 _01151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10162_ _02403_ _02421_ _02416_ _02422_ _02423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_TAPCELL_ROW_7_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09138__A1 _01270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14131__A1 _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10143__I _01555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14970_ _06940_ _06941_ _06942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10093_ _01070_ _02356_ _02357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09689__A2 _02071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13921_ _04272_ _05208_ _05923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08992__S0 _01149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16640_ channels.lfsr\[0\]\[22\] _08390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_92_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08548__I clk_trg\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13852_ _03284_ _05853_ _05854_ _05855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_92_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15631__A1 _02029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12803_ _04723_ _04726_ _04809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_16571_ _08342_ _08348_ _08301_ _08350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13783_ _05700_ _05786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_54_clk clknet_5_10__leaf_clk clknet_leaf_54_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10995_ _03219_ _03220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15522_ _07452_ _07463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_12734_ _04739_ _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_96_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15453_ _07386_ _07390_ _07399_ _07400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_61_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12665_ _04657_ _04659_ _04655_ _04671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XPHY_EDGE_ROW_106_Left_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_155_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12748__A2 _04753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14404_ _05975_ _06401_ _06402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11616_ _03662_ _03712_ _03716_ _00431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15384_ _07315_ _07329_ _07336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_108_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09613__A2 _01937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12596_ _04297_ _04599_ _04601_ _04353_ _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_136_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17123_ _00193_ clknet_leaf_119_clk channels.pw2\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_14335_ _06332_ _05570_ _06225_ _06333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11547_ _03657_ _03669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17054_ _00124_ clknet_leaf_212_clk channels.lfsr\[1\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14266_ _06263_ _06264_ _06265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_11478_ _03612_ _01571_ _03622_ _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16005_ _07799_ _07794_ _07885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13217_ _05219_ _05221_ _05218_ _05223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10429_ _02689_ _02680_ _02690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_59_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14197_ _06122_ _06134_ _06196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11184__A1 _03394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13148_ _05122_ _05125_ _05153_ _05154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_115_Left_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10931__A1 channels.sample1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13079_ _05063_ _05083_ _05085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16907_ channels.exp_counter\[3\]\[2\] _00983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15065__B _06899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16838_ _00928_ _03731_ tt_um_rejunity_sn76489.clk_counter\[1\] _00930_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16769_ _03491_ net12 _00882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16675__I _06978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_45_clk clknet_5_2__leaf_clk clknet_leaf_45_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09310_ _01620_ _01729_ _01731_ _01623_ _00106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_76_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09241_ channels.lfsr\[0\]\[13\] _01676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_111_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09172_ channels.lfsr\[0\]\[3\] _01617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13936__A1 _04446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_155_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13539__I _05543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput18 net18 DAC_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_12_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12443__I _04372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput29 net29 bus_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14113__A1 _04711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08956_ _01254_ _01421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08887_ _01356_ _01357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09540__A1 _01919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09508_ _01898_ _01899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_79_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_175_3624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_175_3635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10780_ _03033_ _03034_ _03035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09439_ _01829_ _01830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_23_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12450_ _04370_ _04454_ _04455_ _04456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_152_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11401_ _02357_ _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_12381_ _04229_ _04386_ _04387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_117_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09927__I _01813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14120_ _06118_ _06119_ _06120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11332_ _03513_ _03522_ _03527_ _00336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_104_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13155__A2 _04315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14051_ _06049_ _06050_ _06051_ _06052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_24_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11263_ _03472_ _03473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13002_ _04462_ _05006_ _05007_ _05008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10214_ _02459_ _02469_ _02474_ _02475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11194_ _03391_ _03392_ _03393_ _03408_ _00317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_30_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10913__A1 channels.sample2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10145_ _02389_ _02405_ channels.pw3\[9\] _02406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_100_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15852__A1 _03735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_54_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17741_ _00811_ clknet_leaf_62_clk tt_um_rejunity_sn76489.control_tone_freq\[0\]\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10076_ filters.cutoff_lut\[15\] _02341_ _02342_ _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14953_ _05647_ _06924_ _06925_ _06926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_89_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13904_ _05821_ _05822_ _05906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17672_ _00742_ clknet_leaf_59_clk tt_um_rejunity_sn76489.tone\[2\].gen.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09531__B2 channels.ctrl_reg3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14884_ filters.low\[27\] _06520_ _03474_ _06863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15604__A1 _01977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16623_ _01650_ _08384_ _08385_ _01653_ _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_13835_ _05836_ _05837_ _05838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_27_clk clknet_5_1__leaf_clk clknet_leaf_27_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16554_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[1\] _08327_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[1\]
+ _08335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13766_ _05767_ _05768_ _05769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_43_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10978_ _03182_ _03203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_70_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15505_ _07446_ _07447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12717_ _04720_ _04721_ _04722_ _04723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_16485_ _08261_ _08275_ _08276_ _08277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_57_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13697_ _05693_ _05696_ _05700_ _05701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_73_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15436_ filters.low\[26\] _06852_ _07384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_66_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12648_ _04354_ _04601_ _04654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15367_ _07299_ _07316_ _07317_ _07277_ _07320_ _07321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_124_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12579_ _04583_ _04584_ _04585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_96_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17106_ _00176_ clknet_leaf_109_clk channels.atk_dec1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_40_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14318_ _06204_ _06209_ _06315_ _06316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_68_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15298_ _07256_ _07257_ _07258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_111_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17037_ _00107_ clknet_leaf_219_clk channels.lfsr\[1\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13146__A2 _05147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_123_Left_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_14249_ _06242_ _06247_ _06248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_81_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13697__A3 _05700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13941__I1 filters.band\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09770__A1 _02112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08810_ channels.ctrl_reg2\[1\] channels.sync_outs\[0\] _01282_ _01283_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09790_ _02105_ _02142_ _02144_ _00177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_175_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08741_ _01222_ _01223_ _01224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09522__A1 channels.atk_dec2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09522__B2 channels.pw3\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08672_ _01155_ _01156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_178_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_178_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_132_Left_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11880__A2 _03964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14949__A3 channels.sample1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_18_clk clknet_5_6__leaf_clk clknet_leaf_18_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__13082__A1 _05080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11342__I _02710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_153_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13909__A1 _04406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09224_ channels.lfsr\[3\]\[10\] _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_170_3532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_170_3543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14582__A1 _05909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09155_ channels.lfsr\[1\]\[1\] _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_130_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_141_Left_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_131_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09086_ _01321_ _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_131_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11148__A1 _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11699__A2 _03789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_168_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11718__S _03784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09988_ _02274_ _02283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_157_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08939_ _01403_ _01404_ _01405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_129_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_150_Right_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_129_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11950_ _04019_ _04028_ _04029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_150_Left_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11320__A1 _03515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10901_ _02365_ _03147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_93_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11881_ _03542_ _03752_ _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13620_ _05145_ _05625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_67_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10832_ _03083_ _03084_ _03085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_156_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13551_ _05494_ _05524_ _05556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_94_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10763_ _03015_ _03017_ _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12502_ _04293_ _04504_ _04182_ _04505_ _04508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_16270_ filters.sample_buff\[11\] _08125_ _08130_ spi_dac_i.spi_dat_buff_0\[7\] spi_dac_i.spi_dat_buff_0\[8\]
+ _08127_ _08132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_66_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13482_ _04480_ _05487_ _05488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10694_ _02907_ _02912_ _02950_ _02951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_81_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15221_ _01762_ channels.sample2\[10\] _07184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14573__A1 _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12433_ net33 _04412_ _04439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_120_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15152_ _07113_ _07117_ _07118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12364_ _04367_ _04369_ _04370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14103_ _06022_ _06056_ _06102_ _06103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_39_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11315_ _03513_ _03508_ _03514_ _00332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_15083_ _07040_ _07050_ _07051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12295_ _04269_ _04301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_56_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14034_ _06033_ _06034_ _06035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_120_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11246_ _03456_ _03225_ _03457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13907__I _05229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09752__A1 _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12351__A3 _04283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11177_ _03244_ _03392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_38_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10128_ _01248_ _02389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15985_ _07840_ _07865_ _07866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_98_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10331__I _02507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17724_ _00794_ clknet_leaf_59_clk tt_um_rejunity_sn76489.control_tone_freq\[2\]\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10059_ _02333_ _02334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14936_ _06909_ _06910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_89_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10114__A2 channels.ring_outs\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17655_ _00725_ clknet_leaf_52_clk tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14867_ _06845_ _06847_ _06848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__16250__A1 _07923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16606_ _08377_ _08378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13818_ _04451_ _05516_ _05821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17586_ _00656_ clknet_leaf_45_clk spi_dac_i.spi_dat_buff_1\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08736__I _01219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14798_ filters.band\[18\] _06785_ _06763_ _06786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16537_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[3\] tt_um_rejunity_sn76489.tone\[1\].gen.counter\[2\]
+ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[1\] tt_um_rejunity_sn76489.tone\[1\].gen.counter\[0\]
+ _08320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_128_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13749_ _03268_ _03375_ _05753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11162__I _03377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16468_ _08257_ _08261_ _08262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_143_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09115__S0 _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13367__A2 _05372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15419_ _07312_ _07367_ _07368_ _00582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_182_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16399_ _08194_ _08211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_182_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11378__A1 _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10050__A1 channels.sus_rel3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12207__B _04212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13119__A2 _05124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09991__A1 _02234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09911_ _02179_ _02227_ _02229_ _00213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09842_ _02180_ _02181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_95_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09773_ _02131_ _02125_ _02132_ _00172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_146_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08724_ channels.exp_periods\[2\]\[1\] _01208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08655_ _01138_ _01139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_139_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_124_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13055__A1 _04900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08586_ _01042_ _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_117_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12168__I _04173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12802__A1 _04792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08482__A1 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09207_ channels.lfsr\[0\]\[8\] _01647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09138_ _01270_ _01537_ _01542_ _01586_ _01587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_121_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09982__A1 _02250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09069_ _01517_ _01518_ _01524_ _01525_ _00071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_11100_ _03318_ _03319_ _03320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12080_ channels.env_counter\[0\]\[8\] _04120_ _04121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11031_ _03254_ _03255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11541__A1 channels.freq2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15770_ _07675_ _07676_ _00625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12982_ _04814_ _04870_ _04872_ _04988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__09940__I _02184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13833__A3 _05145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14721_ filters.band\[12\] _05540_ _05541_ _06715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11933_ _03879_ _03874_ _04015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_59_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17440_ _00510_ clknet_leaf_153_clk channels.accum\[3\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14652_ filters.band\[31\] _04634_ _06647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11864_ _03950_ _03951_ _03952_ _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13603_ _05479_ _05480_ _05608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_157_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12078__I _04103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17371_ _00441_ clknet_leaf_209_clk channels.env_vol\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10815_ _03067_ _03068_ _03069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16773__I _00884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14583_ _04806_ _05448_ _06579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11795_ _01149_ _03886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_28_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16322_ _08159_ _08160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_138_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13534_ _04159_ _05540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10746_ _02676_ _02872_ _03002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16535__A2 _08315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16253_ _07923_ _08120_ _00664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13349__A2 _05354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13465_ _04451_ _04405_ _05471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10677_ _02931_ _02934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09387__I net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08505__B _01032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15204_ _07165_ _07166_ _07167_ _07168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_93_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12416_ _04343_ _04344_ _04422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_93_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16184_ _07761_ _07875_ _07878_ _08058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_51_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13396_ _05399_ _05400_ _05402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_152_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15135_ _07069_ _07099_ _07100_ _07101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_12347_ _04313_ _04353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_142_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15066_ _07032_ _07034_ _00563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12278_ _04252_ _04264_ _04283_ _04284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_71_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15510__A3 _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14017_ _06015_ _06016_ _06017_ _06018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_11229_ _03440_ _03224_ _03441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_156_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15968_ _07783_ _07805_ _07849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_164_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_4_clk_I clknet_5_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10099__A1 _02359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17707_ _00777_ clknet_leaf_229_clk channels.lfsr\[0\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14919_ _06894_ _06885_ _06895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_37_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15899_ _07776_ _07779_ _07780_ _07781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__11835__A2 _03925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17638_ _00708_ clknet_5_19__leaf_clk channels.ch3_env\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__13037__A1 _04992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_172_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13588__A2 _04850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17569_ _00639_ clknet_leaf_34_clk filters.low\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_102_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16526__A2 _08263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09964__A1 channels.pw3\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08767__A2 _01090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_148_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_165_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11523__A1 channels.pw1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10326__A2 _02385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09825_ channels.freq2\[11\] _02164_ _02167_ _02169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15762__I _07332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16462__A1 _08136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15265__A2 _02056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09756_ channels.ctrl_reg1\[6\] _02117_ _02120_ _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09760__I _01780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08707_ channels.exp_counter\[0\]\[4\] channels.exp_counter\[1\]\[4\] channels.exp_counter\[2\]\[4\]
+ channels.exp_counter\[3\]\[4\] _01175_ _01172_ _01191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_119_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09687_ _02065_ _02070_ _02071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15017__A2 filters.filt_1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08638_ channels.env_vol\[3\]\[0\] _01130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_90_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08569_ _01085_ _01086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_166_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10600_ _02641_ _02775_ _02859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11580_ _03673_ _03687_ _03692_ _00419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_36_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10531_ _02686_ _02624_ _02765_ _02791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_49_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12626__I _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13250_ _05186_ _05256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10462_ _02685_ _02703_ _02600_ _02708_ _02723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__13200__A1 _05142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12201_ filters.res_lut\[2\] _04169_ _04207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09955__A1 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13181_ _05186_ _05187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_33_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10393_ _02599_ _02628_ _02642_ _02654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_12132_ channels.accum\[3\]\[14\] _04148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09707__A1 channels.freq1\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12361__I _04366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12063_ _04017_ _04105_ _04110_ _00484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16940_ _00019_ clknet_leaf_220_clk channels.lfsr\[3\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11514__A1 _03511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11014_ _03238_ _03239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_159_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16871_ _01180_ _00938_ _00958_ _00837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15256__A2 _07216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_240_clk clknet_5_18__leaf_clk clknet_leaf_240_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15822_ _06905_ _07640_ _07712_ _00641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_5_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15605__C _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15753_ _06608_ _07664_ _07665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12965_ _04619_ _04966_ _04969_ _04971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_87_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11916_ _03855_ _03998_ _03999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14704_ _06602_ _06697_ _06692_ _06698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_15684_ _07603_ _07609_ _07611_ _07613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_12896_ _03332_ _04371_ net60 _04902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_158_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17423_ _00493_ clknet_leaf_149_clk channels.env_counter\[0\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14635_ _05624_ _05281_ _06630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_47_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11847_ _03744_ _03937_ _03938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_64_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17354_ _00424_ clknet_leaf_96_clk channels.pw3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14566_ _06432_ _06445_ _06562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_64_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11778_ _03801_ _03868_ _03869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12242__A2 _04245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16305_ channels.env_counter\[3\]\[8\] _08150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_126_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13517_ _05499_ _05522_ _05523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_126_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11450__B1 _01448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10729_ _02951_ _02968_ _02985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_67_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17285_ _00355_ clknet_leaf_162_clk channels.accum\[2\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13990__A2 _05990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14497_ _06490_ _06493_ _06494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_153_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16236_ _08101_ _08106_ _08107_ _08108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_42_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13448_ _05445_ _05453_ _05454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_180_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10005__A1 _02245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16167_ _08038_ _08039_ _08041_ _08042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10056__I _02330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13379_ _05384_ _05385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14790__I1 filters.band\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15118_ _07083_ _07084_ _07085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_142_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16098_ _07969_ _07972_ _07975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15049_ _01769_ channels.sample3\[4\] _07018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09066__B _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_78_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09610_ _01892_ _01997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_231_clk clknet_5_20__leaf_clk clknet_leaf_231_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_143_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_160_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_160_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09541_ _01823_ _01930_ _00142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_92_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09472_ channels.sus_rel3\[0\] _01859_ _01862_ channels.pw2\[8\] _01863_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_149_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_121_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09634__B1 _01970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08988__A2 _01443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12446__I _04451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14930__A1 _06769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10547__A2 _02590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12181__I _04186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13497__A1 _04295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_180_3715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_1168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_180_3726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09808_ _01813_ _02157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_222_clk clknet_5_20__leaf_clk clknet_leaf_222_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_210_clk_I clknet_5_20__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09739_ _02105_ _02107_ _02109_ _00161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_2_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13941__S _05179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12750_ _04741_ _04743_ _04756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_9_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12472__A2 _04476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11701_ channels.atk_dec3\[4\] _01078_ _03780_ channels.atk_dec2\[4\] _01291_ channels.atk_dec1\[4\]
+ _03792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA_clkbuf_leaf_225_clk_I clknet_5_20__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14749__A1 _03468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_178_3688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12681_ _04589_ _04590_ _04686_ _04687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14836__I _06760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_15__f_clk_I clknet_3_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14420_ _06325_ _06329_ _06416_ _06417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_49_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11632_ _03677_ _03719_ _03726_ _00437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_154_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13421__A1 _05405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14351_ _06240_ _06248_ _06349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11563_ _03679_ _03681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_80_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11983__A1 _04044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13302_ _04384_ _04816_ _05308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17070_ _00140_ clknet_leaf_99_clk filters.mode_vol\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10514_ _02768_ _02769_ _02773_ _02774_ _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_14282_ _06280_ _06281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_11494_ _03624_ _03632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_21_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16021_ _07849_ _07862_ _07901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15667__I _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09928__A1 channels.sus_rel2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13233_ _05235_ _05238_ _05239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14921__A1 _06722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10445_ _01162_ _02559_ _02705_ _02706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13164_ _05121_ _05126_ _05170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10376_ _02529_ _02634_ _02636_ _02637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_103_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16674__A1 _08356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12115_ _04139_ _00507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13095_ _05099_ _04906_ _05100_ _05101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16923_ _00971_ channels.exp_periods\[0\]\[4\] _00986_ _00992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12046_ channels.adsr_state\[3\]\[0\] _04099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_88_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_213_clk clknet_5_21__leaf_clk clknet_leaf_213_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_16854_ _03096_ _02752_ _00942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_46_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15805_ _06848_ _07690_ _07702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16785_ _08441_ _08442_ _00880_ _00893_ _00881_ _00894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_13997_ _05905_ _05935_ _05998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_66_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12948_ _04493_ _04954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_66_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15736_ _07636_ _07652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13660__A1 _04645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15667_ _03940_ _07597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12879_ _03253_ _04224_ _04884_ _04885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_157_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15401__A2 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17406_ _00476_ clknet_leaf_130_clk channels.env_counter\[1\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14618_ _06517_ _06596_ _06612_ _06613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_15598_ _07532_ _07533_ _07534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17337_ _00407_ clknet_leaf_103_clk channels.freq2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14549_ filters.band\[30\] _04506_ _06545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10777__A2 _02777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17268_ _00338_ clknet_leaf_153_clk channels.adsr_state\[0\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16219_ _08088_ _08091_ _08092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_114_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12518__A3 _04296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17199_ _00269_ clknet_leaf_168_clk channels.sync_outs\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11726__A1 channels.atk_dec3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09575__I _01943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11726__B2 channels.atk_dec2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_1168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15468__A2 _07030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08972_ channels.accum\[0\]\[10\] _01435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13825__I _05469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_204_clk clknet_5_22__leaf_clk clknet_leaf_204_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_120_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11337__S0 _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09524_ channels.freq1\[1\] _01855_ _01857_ channels.ctrl_reg1\[1\] _01914_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12454__A2 _04458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13651__A1 _05553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09455_ _01786_ net1 _01845_ _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_19_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08654__I _00009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09386_ net4 _01784_ _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_19_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09083__A1 _01323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_173_3596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11965__A1 _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16804__C _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15156__A1 _05379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_91_clk_I clknet_5_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13706__A2 _05621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14903__A1 _06614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_18_Left_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_134_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11717__A1 _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10230_ _02461_ _02462_ _02491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_14_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11812__S1 _03842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16656__A1 _08356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10161_ _02360_ _02394_ _02413_ _01553_ _02422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_7_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10940__A2 _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11964__B _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10092_ _01082_ _02356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_96_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13920_ _05835_ _05838_ _05921_ _05922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_96_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08897__B2 channels.freq1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13851_ _03282_ _03220_ _05854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08992__S1 _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_27_Left_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12802_ _04792_ _04807_ _04808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_clkbuf_leaf_164_clk_I clknet_5_28__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16570_ _08342_ _08348_ _08349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13782_ _05703_ _05783_ _05784_ _05785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10994_ _03218_ _03219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_57_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15521_ filters.sample_buff\[0\] _07458_ _07462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_84_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12733_ filters.high\[13\] filters.band\[13\] _04710_ _04739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_44_clk_I clknet_5_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15452_ _07373_ _06767_ _07384_ _07399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_26_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12664_ _04647_ _04651_ _04664_ _04669_ _04670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__15395__A1 _07062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14403_ _06298_ _06400_ _06401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_179_clk_I clknet_5_18__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11615_ channels.pw2\[1\] _03713_ _03714_ _03716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_182_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09074__A1 _01323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15383_ filters.high\[22\] _06919_ _07335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12595_ _04600_ _04601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_182_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10759__A2 _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17122_ _00192_ clknet_leaf_116_clk channels.freq2\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA_clkbuf_leaf_59_clk_I clknet_5_8__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14334_ _04355_ _06332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_182_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11546_ _02149_ _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_128_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17053_ _00123_ clknet_leaf_231_clk channels.lfsr\[1\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_102_clk_I clknet_5_13__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14265_ _04644_ _06261_ _06264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_151_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11477_ channels.accum\[1\]\[23\] _03590_ _03622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14007__S _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16004_ _07881_ _07883_ _07884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13216_ _05218_ _05219_ _05221_ _05222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_10428_ _02675_ _02679_ _02689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_164_Right_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_14196_ _06107_ _06121_ _06195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_59_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12381__A1 _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11184__A2 _03395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13147_ _05123_ _05124_ _05153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_0_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10359_ _01657_ _02386_ _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_117_clk_I clknet_5_27__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13078_ _05063_ _05083_ _05084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12029_ _04041_ _04084_ _04089_ _00471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_139_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16906_ _00982_ _00848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_164_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16837_ _00928_ _03732_ _00929_ _00832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_75_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15860__I _07742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16768_ _01811_ net15 _00881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13633__A1 _05604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_88_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15719_ _07639_ _07640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16699_ _08434_ _08438_ _08439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_180_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09240_ channels.lfsr\[2\]\[14\] _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_173_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_155_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09171_ channels.lfsr\[2\]\[4\] _01616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13936__A2 _04766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_116_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_151_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput19 net19 DAC_dat_1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_113_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_131_Right_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_101_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16638__A1 _01710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08955_ _01337_ _01418_ _01419_ _01420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__13555__I _04645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08886_ _01354_ _01355_ _01356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__13872__A1 _05846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09540__A2 _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10150__A3 channels.pw3\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09507_ _01856_ _01860_ _01898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_3625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_3636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09438_ _01825_ _01826_ _01828_ _01829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_82_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_136_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13927__A2 _05229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09369_ _01769_ _01770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11400_ _03577_ _03569_ _01503_ _03570_ _00354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_145_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12380_ _04385_ _04386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_34_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11331_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[2\] _03523_ _03517_ _03527_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10610__A1 _01556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14050_ _04325_ _05947_ _06051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13155__A3 _04271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11262_ _03471_ _03472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_30_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13001_ _04979_ _04978_ _05007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_162_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10213_ _01509_ _02473_ _02458_ _01498_ _02474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_28_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11193_ _03404_ _03407_ _03408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09943__I _02187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10144_ _01272_ _02405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14104__A2 _06041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17740_ _00810_ clknet_leaf_54_clk tt_um_rejunity_sn76489.control_tone_freq\[0\]\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10075_ _02324_ _02340_ _02344_ _00262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14952_ _01768_ channels.sample3\[0\] _06925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13903_ _05825_ _05842_ _05904_ _05905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_17671_ _00741_ clknet_leaf_79_clk tt_um_rejunity_sn76489.tone\[2\].gen.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14883_ _06706_ _06862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_159_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_30__f_clk_I clknet_3_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16622_ _01645_ _08384_ _08385_ _01647_ _00768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_13834_ _03363_ _04854_ _05731_ _05837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_138_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13615__A1 _03364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16553_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[2\] _08327_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[2\]
+ _08334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13765_ _05563_ _05663_ _05675_ _05768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_130_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10977_ _03191_ _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09295__A1 _01282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15504_ _07443_ _07444_ _07445_ _03729_ _07446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_127_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12716_ _03288_ _04316_ _04197_ _04722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_70_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16484_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[1\] _08268_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[1\]
+ _08276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13696_ _05697_ _05698_ _05699_ _05700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_26_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_155_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15435_ filters.low\[26\] _07383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12647_ _04535_ _04648_ _04653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_25_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15366_ _07307_ _07318_ _07319_ _07320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_12578_ _04540_ _04542_ _04536_ _04584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_25_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17105_ _00175_ clknet_leaf_108_clk channels.atk_dec1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_11529_ channels.pw1\[7\] _03650_ _03652_ _03656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14317_ _06210_ _06214_ _06315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_15297_ _07250_ _07255_ _06982_ _07257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17036_ _00106_ clknet_leaf_221_clk channels.lfsr\[1\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14248_ _06245_ _06246_ _06247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_180_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11788__S0 _01151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14179_ _03330_ _06177_ _06178_ _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_74_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08740_ _01169_ _01206_ _01223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08671_ _01154_ _01155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_75_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13606__A1 _05158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14949__A4 channels.sample2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_157_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09223_ channels.lfsr\[1\]\[10\] _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_153_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13909__A2 _04929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_170_3533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09154_ channels.lfsr\[0\]\[1\] _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_99_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_170_3544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12188__A4 filters.high\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10199__A3 channels.pw2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09085_ _01532_ _01518_ _01539_ _01525_ _00073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_142_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12896__A2 _04371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_168_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09987_ _02274_ _02282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_122_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08938_ _01396_ _01394_ _01402_ _01404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__12648__A2 _04601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_129_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08869_ channels.freq2\[2\] _01275_ _01287_ channels.freq1\[2\] _01340_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_28_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10900_ _02366_ _02880_ _03146_ _00285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11880_ _03960_ _03964_ _03966_ _00445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15433__C _06917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10831_ _03055_ _03056_ _03079_ _03084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13550_ _05442_ _05455_ _05554_ _05555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_137_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10762_ _02979_ _03016_ _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12501_ _04504_ _04206_ _04505_ _04506_ _04507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_66_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09029__A1 _01422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13481_ _04882_ _05487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_137_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10693_ _02899_ _02906_ _02950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_82_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15220_ _01771_ channels.sample3\[10\] _07183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12432_ _04436_ _04427_ _04437_ _04438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_129_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15151_ _07114_ _07078_ _07116_ _07117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_129_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12363_ _04368_ _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_106_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14102_ _06024_ _06055_ _06102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11314_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[2\] _03509_ _03503_ _03514_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14325__A2 _04924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15082_ _07043_ _07049_ _07050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_121_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12294_ _04270_ _04298_ _04299_ _04300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14033_ _04750_ _04884_ _06034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_56_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11245_ filters.band\[14\] _03456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_91_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10898__A1 _02366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11176_ filters.sample_filtered\[10\] _03391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_10127_ _01534_ _02382_ _02387_ _02388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_98_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15984_ _07845_ _07864_ _07865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_17723_ _00793_ clknet_leaf_53_clk tt_um_rejunity_sn76489.chan\[0\].attenuation.in
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11698__I0 channels.atk_dec1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10058_ _01750_ _02333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14935_ _06908_ _06909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_145_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17654_ _00724_ clknet_leaf_64_clk tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15589__A1 channels.sample3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14866_ _06836_ _06846_ _06847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_58_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16605_ _01724_ _08374_ _08377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13817_ _05158_ _05074_ _05820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_17585_ _00655_ clknet_leaf_46_clk spi_dac_i.spi_dat_buff_1\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09268__B2 _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13064__A2 _05069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14797_ _06760_ _06785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11443__I _01104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16536_ _02347_ _08315_ _08319_ _00748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13748_ _05751_ _05752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_174_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16455__B _08252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16467_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[0\] _08260_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[0\]
+ _08261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_14_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13679_ _05591_ _05599_ _05682_ _05683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_26_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15418_ filters.high\[24\] _07310_ _07356_ _07368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09115__S1 _01154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16398_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[6\] _08209_ _08210_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_170_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09440__A1 net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15349_ filters.low\[19\] _06498_ _07304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_76_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15513__A1 _03263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12327__A1 _03302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09910_ channels.sus_rel2\[0\] _02228_ _02224_ _02229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_22_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17019_ _00098_ clknet_leaf_235_clk channels.lfsr\[2\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09841_ _02088_ _01862_ _02180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__13319__B _05324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09772_ channels.atk_dec1\[3\] _02126_ _02129_ _02132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13827__A1 _04864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_146_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08723_ channels.exp_periods\[0\]\[1\] channels.exp_periods\[1\]\[1\] _01187_ _01207_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_179_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08654_ _00009_ _01138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__16241__A2 _07722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08585_ _01100_ _01101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14865__S _03473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13055__A2 _04905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_92_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12802__A2 _04807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_174_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09206_ channels.lfsr\[2\]\[9\] _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_49_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08662__I _01145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09137_ _01585_ _01586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_161_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09068_ _01254_ _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_163_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_13__f_clk clknet_3_3_0_clk clknet_5_13__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11030_ _03253_ _03254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_34_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13818__A1 _04451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12981_ _04983_ _04984_ _04986_ _04987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14720_ net30 _06713_ _06714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11932_ _04008_ _04010_ _04014_ _00449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_169_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14651_ _06644_ _06645_ _06646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11863_ _03749_ _03946_ _03952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_68_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11263__I _03472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13602_ _05470_ _05605_ _05606_ _05607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10814_ _03065_ _03066_ _03068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17370_ _00440_ clknet_leaf_166_clk channels.clk_div\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11794_ _03804_ _03845_ _03885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14582_ _05909_ _05367_ _06578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16321_ _02363_ _03936_ _01821_ _08159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_95_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_165_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10745_ _02657_ _02823_ _03001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13533_ _05537_ _05538_ _05539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_137_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16252_ filters.sample_buff\[5\] _08115_ _08117_ spi_dac_i.spi_dat_buff_0\[1\] spi_dac_i.spi_dat_buff_0\[2\]
+ _08119_ _08120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_13464_ _05158_ _05469_ _05470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_168_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15743__A1 _03345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10676_ _02882_ _02932_ _02933_ _00274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_153_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12557__A1 _04468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12415_ _04301_ _04420_ _04421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15203_ _03374_ _07133_ _07167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_93_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16183_ _08033_ _08055_ _08056_ _08057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09422__A1 filters.hp vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13395_ _05399_ _05400_ _05401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_93_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12346_ _04328_ _04348_ _04351_ _04352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_65_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15134_ _07072_ _07076_ _07100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_181_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15065_ filters.high\[5\] _07033_ _06899_ _07034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12277_ _04270_ _04275_ _04282_ _04283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XTAP_TAPCELL_ROW_71_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14016_ _04230_ _05505_ _06017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_71_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11228_ filters.band\[13\] _03440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__09281__S0 _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11159_ _03217_ _03375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_175_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15967_ _07810_ _07816_ _07846_ _07847_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[1\]
+ _07848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_175_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17706_ _00776_ clknet_leaf_235_clk channels.lfsr\[0\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14918_ _06878_ _06894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_78_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15898_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[3\] _07766_ _07780_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_72_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17637_ _00707_ clknet_leaf_208_clk channels.ch3_env\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_59_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14849_ _06795_ _06808_ _06814_ _06825_ _06831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_176_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_86_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17568_ _00638_ clknet_leaf_34_clk filters.low\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15801__C _07269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16519_ _08300_ _08304_ _08306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09661__A1 channels.pw1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17499_ _00569_ clknet_leaf_6_clk filters.high\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09661__B2 channels.ctrl_reg1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15734__A1 _03310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_30_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16913__B _01043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_170_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09964__A2 _02266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_148_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_165_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10252__I _02512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09824_ _02112_ _02163_ _02168_ _00187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__16462__A2 _07924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09755_ _02093_ _02120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_20_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13276__A2 _05281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08706_ _01186_ _01189_ _01190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09686_ _02066_ _02067_ _02068_ _02069_ _02070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08657__I _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15017__A3 channels.sample1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08637_ _01129_ _00035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_68_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12179__I _04184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14225__A1 _04893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08568_ channels.accum\[0\]\[23\] channels.accum\[1\]\[23\] channels.accum\[2\]\[23\]
+ channels.accum\[3\]\[23\] _00009_ _00010_ _01085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_92_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08499_ _01009_ _01021_ _01025_ _01027_ _01028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_153_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10530_ _02738_ _02781_ _02789_ _02790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10461_ _02713_ _02721_ _02716_ _02722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_51_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09404__A1 _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13200__A2 _05147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12200_ _04182_ _04206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13180_ _05185_ _05186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10392_ _02555_ _02503_ _02653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_62_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12131_ _04147_ _00515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_62_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12062_ channels.env_counter\[0\]\[1\] _04108_ _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11013_ _03180_ _03238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_16870_ _00939_ _00957_ _00958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_15821_ filters.low\[31\] _07631_ _07700_ _07712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11278__A1 _02308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08567__I _01083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15752_ _07663_ _07664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12964_ _04619_ _04966_ _04969_ _04970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_73_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14703_ _06400_ _06502_ _06697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11915_ _03992_ _03889_ _03993_ _03997_ _03998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_15683_ _07603_ _07609_ _07611_ _07612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_12895_ _04367_ _04268_ _04901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17422_ _00492_ clknet_leaf_150_clk channels.env_counter\[0\]\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_158_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14634_ _04447_ _05766_ _06629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11846_ _03936_ _03937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_129_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17353_ _00423_ clknet_leaf_96_clk channels.pw3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_64_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11777_ _03794_ _03845_ _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14565_ _06417_ _06431_ _06561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09398__I _01752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16304_ _08149_ _00686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_82_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13516_ _05508_ _05521_ _05522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10728_ _02951_ _02968_ _02984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_17284_ _00354_ clknet_leaf_154_clk channels.accum\[2\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14496_ _06491_ _06492_ _06493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16235_ _08101_ _08106_ _07741_ _08107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_180_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13447_ _05451_ _05452_ _05453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10659_ _02915_ _02916_ _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16166_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[3\] _07776_ _08040_
+ _08041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13378_ _05383_ _05056_ _05384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_106_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13648__I _01822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15117_ _07026_ _07036_ _07060_ _07084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12329_ _03271_ _04253_ _04241_ _04335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_50_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16097_ _07838_ _07973_ _07974_ _00654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_121_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15048_ _06987_ _07016_ _07017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_103_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12702__A1 _04701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16444__A2 _08244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16895__S _00975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13258__A2 _05263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16999_ _00078_ clknet_leaf_189_clk channels.accum\[0\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_160_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09540_ _01919_ _01923_ _01929_ net23 _01909_ _01930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_TAPCELL_ROW_160_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09471_ _01861_ _01862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_149_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14207__A1 _04737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_121_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10492__A2 _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09634__A1 channels.sus_rel3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09634__B2 channels.freq1\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12233__A3 _04238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_178_Right_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11441__A1 _03600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09101__I _01549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10247__I _02507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_119_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_144_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13558__I _04562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12941__A1 _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12462__I _04390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_160_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_180_3716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_3727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09771__I _01776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09807_ _02155_ _02151_ _02156_ _00182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13249__A2 _05254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09738_ channels.ctrl_reg1\[0\] _02108_ _02094_ _02109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09322__B1 _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09873__A1 _02150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09669_ _01934_ net28 _02036_ _02054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_167_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11700_ _03532_ _03791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_178_3678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12680_ _04559_ _04560_ _04586_ _04686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14749__A2 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_178_3689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11631_ channels.pw2\[7\] _03720_ _03722_ _03726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_167_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12637__I _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13421__A2 _05415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_145_Right_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11562_ _03679_ _03680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_119_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14350_ _06242_ _06247_ _06348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10513_ _02499_ _02774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_13301_ _05212_ _05215_ _05306_ _05307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14281_ _06164_ _06167_ _06280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_52_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11493_ _03515_ _03625_ _03631_ _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__16371__A1 channels.ch3_env\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16020_ _07850_ _07852_ _07854_ _07860_ _07900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__09946__I _02174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13232_ _05236_ _05237_ _05238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10444_ _01162_ _02558_ _02705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08850__I _01321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14073__B _05968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13163_ _05121_ _05126_ _05169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12372__I _04377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10375_ _01156_ _02635_ _02636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12114_ channels.accum\[3\]\[5\] _04139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13094_ _04878_ _04891_ _05100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14685__A1 _06675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12045_ _04072_ _04075_ _04098_ _00478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11499__A1 channels.freq1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16922_ _00991_ _00855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_88_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16853_ _02707_ _03742_ _00941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__10171__A1 _01541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15804_ _06841_ _07640_ _07701_ _00634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12448__B1 _04453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16784_ _01805_ net12 _00893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13996_ _05984_ _05996_ _05997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_137_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_66_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15735_ _07650_ _07651_ _00615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_99_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12947_ _04475_ _04482_ _04953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_73_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11671__A1 channels.sus_rel1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15666_ _07586_ _07596_ _07573_ _00601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12878_ _04816_ _04884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_17405_ _00475_ clknet_leaf_149_clk channels.env_counter\[1\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14617_ _06611_ _06595_ _06612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11829_ _03842_ _03916_ _03919_ _03920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_7_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15597_ _07524_ _07521_ _07531_ _07533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_117_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17336_ _00406_ clknet_leaf_100_clk channels.freq2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14548_ _06380_ _04600_ _06544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_172_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09092__A2 _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_112_Right_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17267_ _00337_ clknet_leaf_70_clk tt_um_rejunity_sn76489.control_tone_freq\[1\]\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15165__A2 channels.sample2\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14479_ _06474_ _06475_ _06476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_102_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13176__A1 _05181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16218_ _08058_ _08089_ _08090_ _08091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_140_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17198_ _00268_ clknet_leaf_168_clk channels.sync_outs\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16149_ _08013_ _08024_ _08025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_51_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08971_ _01422_ _01433_ _01434_ _00064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13479__A2 _04884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14428__A1 _06420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13100__A1 filters.cutoff_lut\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11337__S1 _01161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09523_ filters.cutoff_lut\[7\] _01849_ _01851_ filters.cutoff_lut\[10\] _01913_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_116_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12454__A3 _04459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09454_ net6 net5 _01845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_94_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09385_ net3 _01784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_93_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14873__S _03473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_5_7__f_clk_I clknet_3_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12206__A3 _04211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_173_3586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_173_3597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15156__A2 _05403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16353__A1 _02356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_104_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10160_ _01555_ _02419_ _02408_ _02420_ _01550_ _02421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_112_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09218__S0 _01142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09138__A3 _01542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10091_ _01065_ _02351_ _02355_ _02354_ _00267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_22_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_76_Right_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__15008__I _06978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13850_ _03376_ _05853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_92_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12801_ _04322_ _04802_ _04806_ _04313_ _04807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_97_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13781_ _05705_ _05739_ _05784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10993_ _03217_ _03218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_69_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15520_ _07446_ _07461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12732_ _04173_ _04737_ _04738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08845__I _01317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15451_ _07395_ _07396_ _07397_ _07398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_26_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12663_ _04665_ _04666_ _04668_ _04669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_61_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14402_ _06396_ _06399_ _06400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11614_ _03710_ _03712_ _03715_ _00430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_65_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15382_ _07331_ _07334_ _00579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_154_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12594_ _04296_ _04600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17121_ _00191_ clknet_leaf_116_clk channels.freq2\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_65_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_85_Right_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_108_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14333_ _06316_ _06330_ _06331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11545_ _03666_ _03658_ _03667_ _00409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_131_clk clknet_5_31__leaf_clk clknet_leaf_131_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_151_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17052_ _00122_ clknet_leaf_232_clk channels.lfsr\[1\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14264_ _06260_ _06262_ _06263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11476_ _01563_ _03615_ _01568_ _03616_ _00386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_16003_ _07792_ _07882_ _07883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11708__A2 _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10427_ _02685_ _02514_ _02687_ _02679_ _02688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_13215_ _04386_ _05220_ _04791_ _04180_ _05221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_33_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14195_ _06136_ _06159_ _06193_ _06194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_150_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16647__A2 _08263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13146_ _05142_ _05147_ net49 _05152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_57_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10358_ _01534_ _02539_ _02619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_143_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10392__A1 _02555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14658__A1 _06614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17545__D _00615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13077_ _05073_ _05082_ _05083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_57_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10289_ _02371_ _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_57_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13330__A1 _05234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_94_Right_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12028_ channels.env_counter\[1\]\[7\] _04085_ _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16905_ channels.exp_counter\[3\]\[1\] _00982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_139_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11446__I _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16836_ _00928_ _03731_ _00877_ _00929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16767_ tt_um_rejunity_sn76489.latch_control_reg\[0\] _01816_ _00880_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13979_ _05892_ _05980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_87_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10447__A2 _02707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15718_ _07629_ _07639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16698_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[9\] _08437_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[9\]
+ _08438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_15649_ _07580_ _07581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_115_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09170_ _01609_ _01611_ _01615_ _01599_ _00082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_127_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_1_Left_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_155_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17319_ _00389_ clknet_leaf_243_clk filters.res_lut\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_122_clk clknet_5_30__leaf_clk clknet_leaf_122_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_12_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_79_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_102_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11130__B _03347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_224_clk_I clknet_5_20__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__17128__CLK clknet_5_27__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08954_ _01411_ _01404_ _01417_ _01419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13321__A1 _04395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08885_ channels.accum\[0\]\[3\] channels.accum\[1\]\[3\] channels.accum\[2\]\[3\]
+ channels.accum\[3\]\[3\] _01308_ _01160_ _01355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
Xclkbuf_leaf_189_clk clknet_5_22__leaf_clk clknet_leaf_189_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__13872__A2 _05848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_239_clk_I clknet_5_16__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input16_I bus_we vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14821__A1 _06769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09506_ filters.mode_vol\[0\] _01791_ _01896_ channels.pw3\[0\] _01897_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08665__I _01148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_175_3626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_175_3637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09437_ _01827_ _01828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_164_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_136_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09368_ _01768_ _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_113_clk clknet_5_15__leaf_clk clknet_leaf_113_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09299_ _01724_ _01721_ _01725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_145_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11330_ _03511_ _03522_ _03526_ _00335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_104_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11261_ _03470_ _03471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_160_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10212_ _02470_ _01099_ _02471_ _02472_ _02473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_13000_ _04465_ _04495_ _05006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_162_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11192_ filters.sample_filtered\[9\] _03385_ _03406_ _03407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_101_1304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10143_ _01555_ _02404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_37_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15301__A2 _06065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10074_ filters.cutoff_lut\[14\] _02341_ _02342_ _02344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_54_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14951_ _06922_ _06923_ _06924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10126__A1 _01632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13902_ _05827_ _05841_ _05904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17670_ _00740_ clknet_leaf_79_clk tt_um_rejunity_sn76489.tone\[2\].gen.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14882_ _06859_ _06861_ _00552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__15065__A1 filters.high\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16621_ _08382_ _08385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13833_ _03349_ _04191_ _05145_ _05836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_173_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16552_ _08237_ _08333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11626__A1 _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13764_ _04667_ _05766_ _05673_ _05767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_35_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10976_ _03197_ _03201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_168_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15503_ _01748_ _03428_ _03476_ _01762_ _07443_ _03237_ _07445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_12715_ _03271_ _04241_ _04376_ _04721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_16483_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[2\] _08268_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[2\]
+ _08275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15368__A2 _07321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13695_ _04222_ _05280_ _05699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15434_ _01932_ _07382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12646_ _04647_ _04651_ _04652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_182_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_104_clk clknet_5_13__leaf_clk clknet_leaf_104_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_26_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15365_ _07303_ _07304_ _07319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12577_ _04581_ _04582_ _04583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_109_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17104_ _00174_ clknet_leaf_109_clk channels.atk_dec1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_53_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14316_ _06312_ _06313_ _06314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11528_ _02326_ _03649_ _03655_ _00404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10601__A2 _02500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15296_ _07250_ _07255_ _07256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_151_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17035_ _00105_ clknet_leaf_217_clk channels.lfsr\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14247_ _04231_ _05891_ _06246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11459_ _02364_ _03612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_110_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11788__S1 _01167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14178_ _03329_ _05853_ _06178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_111_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13129_ _05103_ _05109_ _05135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_input8_I bus_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08670_ _01153_ _01154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_79_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15056__A1 _04992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_90_clk_I clknet_5_12__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16819_ _02102_ _00919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14487__I filters.band\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13606__A2 _05516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14803__A1 _06769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11617__A1 channels.pw2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_157_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_46_Left_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09222_ channels.lfsr\[0\]\[10\] _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_118_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14031__A2 _04403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09153_ channels.lfsr\[2\]\[2\] _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_170_3534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_170_3545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09084_ _01535_ _01538_ _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_131_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_163_clk_I clknet_5_28__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12345__A2 _04283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_55_Left_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_101_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12470__I _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_168_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09986_ _02215_ _02275_ _02281_ _00236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_178_clk_I clknet_5_18__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08937_ _01396_ _01394_ _01402_ _01403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_129_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08868_ channels.freq3\[2\] _01075_ _01339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_58_clk_I clknet_5_8__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16244__B1 _07728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16795__A1 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_101_clk_I clknet_5_13__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08799_ channels.clk_div\[1\] _01272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_10830_ _03047_ _03082_ _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_168_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_64_Left_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10761_ _03012_ _03016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_94_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12820__A3 _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12500_ _04187_ _04506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_clkbuf_leaf_116_clk_I clknet_5_26__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13480_ _04278_ _05208_ _05486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10692_ _02947_ _02948_ _02949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_180_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12431_ _04328_ _04363_ _04413_ _04437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_152_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15150_ _07115_ _07116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_35_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12362_ _04241_ _03270_ _04368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_62_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14101_ _06089_ _06100_ _06101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_95_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11313_ _02187_ _03513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_39_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12293_ _04281_ _04291_ _04293_ _04296_ _04299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_TAPCELL_ROW_39_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15081_ _07048_ _07049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_73_Left_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_56_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14032_ _06031_ _06032_ _06033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_11244_ filters.low\[14\] _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_121_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15177__B _07086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10347__A1 _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11175_ _03372_ _03327_ _03328_ _03390_ _00316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_38_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10898__A2 _02831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15286__A1 _05968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10126_ _01632_ _02386_ _02387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15825__A3 _03731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15983_ _07848_ _07863_ _07864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__16787__I _00895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17722_ _00792_ clknet_leaf_62_clk tt_um_rejunity_sn76489.tone\[0\].gen.counter\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14884__I1 _06520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10057_ _02330_ _02332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14934_ _06907_ _06908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11847__A1 _03744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17653_ _00723_ clknet_leaf_51_clk tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14865_ filters.low\[25\] filters.band\[25\] _03473_ _06846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_82_Left_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16604_ _08375_ _08376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_159_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13816_ _05720_ _05817_ _05818_ _05819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_17584_ _00654_ clknet_leaf_46_clk spi_dac_i.spi_dat_buff_1\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09268__A2 _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14796_ _06748_ _06783_ _06784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_159_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13064__A3 _04341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16736__B _08459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16535_ _02347_ _08315_ _08318_ _08319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13747_ _05750_ _05751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10959_ _03180_ _03182_ _03183_ _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_85_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16466_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[9\] tt_um_rejunity_sn76489.tone\[2\].gen.counter\[8\]
+ _08258_ _08259_ _08260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_45_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13678_ _05594_ _05598_ _05682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_171_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15417_ _07362_ _07366_ _07367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__12555__I _04500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12629_ _03256_ _04566_ _04633_ _04634_ _04635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
X_16397_ _08197_ _08209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_143_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15348_ filters.low\[18\] _06396_ _07303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09440__A2 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_170_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16471__B _07740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_91_Left_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14770__I _04159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15279_ _07029_ _07240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_110_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17018_ _00097_ clknet_leaf_231_clk channels.lfsr\[2\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12327__A2 _04332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09840_ _02104_ _02179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12290__I _04295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08951__A1 _01414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09771_ _01776_ _02131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13827__A2 _05721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08722_ channels.exp_counter\[0\]\[1\] channels.exp_counter\[1\]\[1\] channels.exp_counter\[2\]\[1\]
+ channels.exp_counter\[3\]\[1\] _01152_ _01168_ _01206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__11838__A1 _01584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08653_ _01137_ _00043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_152_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_124_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08584_ _01095_ _01099_ _01100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_117_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09104__I _01555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14945__I _01932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09205_ _01639_ _01634_ _01645_ _01627_ _00087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_63_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09136_ _01584_ _01585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_32_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17466__CLK clknet_5_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09067_ _01436_ _01522_ _01523_ _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_60_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13515__A1 _05514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09969_ _02252_ _02265_ _02269_ _00231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13818__A2 _05516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11829__A1 _03842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12980_ _04980_ _04985_ _04982_ _04986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11931_ channels.env_counter\[2\]\[0\] _04013_ _04014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_1230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14650_ _06549_ _06557_ _06645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11862_ _03945_ _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13601_ _05471_ _05472_ _05606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_0_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10813_ _03065_ _03066_ _03067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_68_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14581_ _04802_ _05501_ _06577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11793_ _03848_ _03884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16320_ _08157_ _08158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_83_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13532_ _05535_ _05536_ _05533_ _05538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10744_ _02710_ _02923_ _03000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09670__A2 _02053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16251_ _07727_ _08119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12006__A1 _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13463_ _04737_ _05469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13203__B1 _05208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10675_ channels.sample3\[3\] _02784_ _02933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15202_ _07134_ _07166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_12414_ _04287_ _04420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12557__A2 _04562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16182_ _08036_ _08052_ _08056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_93_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13394_ _05132_ _05192_ _05194_ _05400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_93_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15133_ _07072_ _07076_ _07099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12345_ _04349_ _04283_ _04350_ _04351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_51_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15064_ _06982_ _07033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_121_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12276_ _04281_ _04201_ _04282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_71_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14015_ _04259_ _05351_ _06016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_71_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11227_ filters.low\[13\] _03439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09281__S1 _01680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08933__B2 channels.freq1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11158_ filters.low\[9\] _03374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_175_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10109_ _01266_ channels.ctrl_reg3\[4\] channels.ctrl_reg1\[4\] _01252_ _02370_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_15966_ _07810_ _07815_ _07847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11089_ filters.sample_filtered\[5\] _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_14917_ _06891_ _03477_ _06892_ _06893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_17705_ _00775_ clknet_leaf_235_clk channels.lfsr\[0\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15897_ _07777_ _07769_ _07778_ _07779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_159_Right_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_69_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17636_ _00706_ clknet_leaf_185_clk channels.exp_counter\[0\]\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_69_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14848_ _06829_ _06830_ _00549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_86_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_86_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17567_ _00637_ clknet_leaf_32_clk filters.low\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14765__I _03472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14779_ _06767_ _06768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_58_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09110__A1 _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16518_ _08300_ _08304_ _08305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_85_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17498_ _00568_ clknet_leaf_13_clk filters.high\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_156_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16449_ _08247_ _08248_ _00732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_rebuffer6_I _05423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16931__A1 _01766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_171_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_182_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_111_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_165_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08924__A1 _01389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09823_ channels.freq2\[10\] _02164_ _02167_ _02168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_129_Left_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_182_3780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09754_ _01807_ _02116_ _02119_ _00166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_126_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08705_ channels.exp_periods\[0\]\[2\] channels.exp_periods\[1\]\[2\] channels.exp_periods\[2\]\[2\]
+ channels.exp_periods\[3\]\[2\] _01187_ _01188_ _01189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__11287__A2 _01003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09685_ channels.pw1\[7\] _02003_ _01996_ channels.pw2\[7\] _02069_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_94_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_93_clk clknet_5_7__leaf_clk clknet_leaf_93_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_126_Right_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08636_ channels.lfsr\[3\]\[22\] _01129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15017__A4 channels.sample2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15280__B _07240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08567_ _01083_ _01084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13984__A1 _05940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12787__A2 _04323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_138_Left_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_175_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08498_ _01026_ _01019_ _01027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_92_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10798__A1 channels.sample3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09652__A2 _02035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_107_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_175_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12195__I _04200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10262__A3 _02522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10460_ _01164_ _02520_ _02720_ _02721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_107_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09119_ _01558_ _01566_ _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_165_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10391_ _02566_ _02611_ _02651_ _02652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_60_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12130_ channels.accum\[3\]\[13\] _04147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12061_ _04010_ _04105_ _04109_ _00483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_147_Left_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09009__I _01469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11012_ _03204_ _03215_ _03237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_99_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_159_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15820_ _06891_ _07697_ _07711_ _07710_ _00640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_5_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15751_ _07635_ _07663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_172_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12963_ _04484_ _04967_ _04968_ _04969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__12475__A1 _04220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14702_ _04161_ _06695_ _06696_ _00537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11914_ _03994_ _03995_ _03996_ _03927_ _03997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_15682_ filters.sample_buff\[13\] _07610_ _07611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_12894_ _04897_ _04898_ _04899_ _04900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_87_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17421_ _00491_ clknet_leaf_150_clk channels.env_counter\[0\]\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_169_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14633_ _04318_ _05980_ _06628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11845_ _03779_ _03935_ _03936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_28_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17352_ _00422_ clknet_leaf_96_clk channels.pw3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14564_ _06540_ _06559_ _06560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_56_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11776_ _03865_ _03866_ _03867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_64_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16303_ channels.env_counter\[3\]\[7\] _08149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13515_ _05514_ _05520_ _05521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_17283_ _00353_ clknet_leaf_164_clk channels.accum\[2\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10727_ _02947_ _02948_ _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_126_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16913__A1 _03744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14495_ _06305_ _06389_ _06492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16234_ _08103_ _08105_ _08106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_152_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13446_ _04642_ _05449_ _05452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_180_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10658_ _02859_ _02862_ _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_140_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16165_ _08014_ _07892_ _07856_ _08040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_180_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13377_ _04629_ _05054_ _05383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10589_ _02750_ _02805_ _02847_ _02713_ _02848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_140_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15116_ _07055_ _07059_ _07083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12328_ _04262_ _04333_ _04334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16096_ spi_dac_i.spi_dat_buff_1\[3\] _07867_ _07921_ spi_dac_i.spi_dat_buff_1\[4\]
+ _07871_ _07974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__14152__A1 _04258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15047_ _06989_ _06990_ _07016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12259_ _04174_ _04265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_43_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_143_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16998_ _00077_ clknet_leaf_156_clk channels.accum\[0\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_160_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11269__A2 _03236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15949_ _07811_ _07816_ _07830_ _07831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__12466__B2 _04471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_75_clk clknet_5_14__leaf_clk clknet_leaf_75_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09331__A1 _01705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09470_ _01785_ _01860_ _01861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_121_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14207__A2 _05731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_121_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17619_ _00689_ clknet_leaf_145_clk channels.env_counter\[3\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_175_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_93_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15955__A2 _07728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13966__A1 _05877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11133__B _03350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13718__A1 _03383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14766__I0 filters.low\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_119_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14391__A1 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer19_I _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12941__A2 _04946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10952__A1 channels.sample1\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14143__A1 _04529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_1197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_180_3717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_3728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09806_ channels.sus_rel1\[5\] _02152_ _02146_ _02156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_157_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08668__I _01151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10180__A2 channels.pw2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15643__A1 channels.sample3\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09737_ _02106_ _02108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_2_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_66_clk clknet_5_11__leaf_clk clknet_leaf_66_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09322__A1 _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09668_ _02047_ _02052_ _02053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_69_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_173_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08619_ _01120_ _00026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12209__A1 _03239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_178_3679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09599_ _01909_ net25 _01986_ _01987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11630_ _03675_ _03719_ _03725_ _00436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13957__A1 _05905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09181__S0 _01605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11561_ _03640_ _01871_ _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_9_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12854__S _04710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13709__A1 _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13300_ _05213_ _05214_ _05306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_42_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10512_ _01550_ _02770_ _02772_ _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_14280_ _06168_ _06279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_11492_ channels.freq1\[3\] _03626_ _03627_ _03631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_150_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13231_ _03382_ _04371_ _04342_ _05237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_10443_ _02684_ _02630_ _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13162_ _05073_ _05082_ _05167_ _05168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10374_ channels.env_vol\[0\]\[7\] channels.env_vol\[1\]\[7\] _02518_ _02635_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_21_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10943__A1 channels.sample1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12113_ _04138_ _00506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_5_24__f_clk_I clknet_3_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10173__I channels.pw1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13093_ _04878_ _04891_ _05099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12044_ channels.env_counter\[1\]\[14\] _04078_ _04098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16921_ _00969_ channels.exp_periods\[0\]\[3\] _00987_ _00991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_137_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09561__A1 channels.pw1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09561__B2 channels.freq2\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10901__I _02365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16852_ _01583_ _03737_ _01092_ _01069_ _00940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__14437__A2 _05671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15634__A1 channels.sample1\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15803_ _07363_ _07631_ _07700_ _07701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16783_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[0\] _00892_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_137_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13995_ _05987_ _05995_ _05996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xclkbuf_leaf_57_clk clknet_5_3__leaf_clk clknet_leaf_57_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15734_ _03310_ _07643_ _07644_ _07651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12946_ _04775_ _04874_ _04951_ _04952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_0_88_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15665_ _07450_ _07594_ _07595_ _07596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12877_ _03199_ _04215_ _04882_ _04883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_75_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17404_ _00474_ clknet_leaf_148_clk channels.env_counter\[1\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14616_ _06519_ _06611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_11828_ _01151_ _03917_ _03918_ _01170_ _03919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_56_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15596_ _07524_ _07521_ _07531_ _07532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_68_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09202__I _01604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17335_ _00405_ clknet_leaf_97_clk channels.pw1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14547_ filters.band\[29\] _05446_ _06543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11759_ _03801_ _03850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17266_ _00336_ clknet_leaf_70_clk tt_um_rejunity_sn76489.control_tone_freq\[1\]\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_102_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14478_ _05982_ _06383_ _06382_ _06475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_154_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13659__I _05570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16217_ _08059_ _08068_ _08090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_24_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13429_ _05360_ _05433_ _05434_ _05435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__13176__A2 _04537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17197_ _00267_ clknet_leaf_79_clk clk_trg\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_102_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11187__A1 filters.high\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16148_ _08017_ _08021_ _08023_ _08024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_80_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_114_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16079_ _07811_ _07906_ _07957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08970_ channels.accum\[0\]\[9\] _01360_ _01434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15095__B _06775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput1 addr[0] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_78_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_48_clk clknet_5_10__leaf_clk clknet_leaf_48_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09522_ channels.atk_dec2\[1\] _01838_ _01842_ channels.pw3\[9\] _01912_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_78_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09453_ _01002_ _01844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_176_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13939__A1 _04176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09384_ _01782_ net5 _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_4_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09607__A2 _01989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10217__A3 channels.pw2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_138_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_173_3587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_149_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08910__S0 _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_173_3598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16353__A2 _03936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10207__B _01481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14116__A1 _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09218__S1 _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10090_ net9 _02351_ _02355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_96_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11350__A1 _02847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15616__A1 channels.sample3\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_39_clk clknet_5_3__leaf_clk clknet_leaf_39_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12800_ _04805_ _04806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13780_ _05705_ _05739_ _05783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10992_ _03188_ _03217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12731_ _04711_ _04737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_69_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11552__I _02154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15450_ _07383_ _06734_ _07397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12662_ _04667_ _04635_ _04646_ _04668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_182_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09022__I _01481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_61_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14401_ _03361_ _06397_ _06398_ _06399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_11613_ channels.pw2\[0\] _03713_ _03714_ _03715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15381_ filters.high\[21\] _07033_ _07333_ _07334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_108_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12593_ _04506_ _04599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_0_clk_I clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17120_ _00190_ clknet_leaf_115_clk channels.freq2\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_14332_ _06325_ _06329_ _06330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_52_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11544_ channels.freq2\[3\] _03659_ _03660_ _03667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_135_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17051_ _00121_ clknet_leaf_230_clk channels.lfsr\[1\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13158__A2 _05157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14263_ _04616_ _06261_ _06146_ _06262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_151_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11475_ _03612_ _01559_ _03621_ _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_162_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16002_ _07788_ _07793_ _07882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_111_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13214_ _04780_ _05220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_150_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10426_ _02686_ _02687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_14194_ _06105_ _06135_ _06193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__10916__A1 channels.sample2\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14812__B _06734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09782__A1 channels.atk_dec1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13145_ _05148_ _05149_ _05150_ _05151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_10357_ _02616_ _02617_ _02618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10392__A2 _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14658__A2 _05982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13076_ _05076_ _05080_ _05081_ _05082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_10288_ _01521_ _02377_ _02549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_100_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09534__A1 channels.pw1\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09534__B2 channels.freq2\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12027_ _04037_ _04084_ _04088_ _00470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16904_ _00981_ _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15607__A1 channels.sample1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16739__B _08459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16835_ tt_um_rejunity_sn76489.clk_counter\[0\] _00928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16280__A1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16766_ _03494_ _00879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13978_ _05899_ _05960_ _05978_ _05979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_87_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12929_ _04876_ _04934_ _04935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_15717_ _05651_ _07637_ _07638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16697_ _08242_ _08400_ _08437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_48_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15648_ filters.sample_buff\[10\] _07579_ _07580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_28_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15579_ channels.sample2\[5\] _03378_ _07515_ _03231_ _07516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_29_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_155_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09065__A3 _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17318_ _00388_ clknet_leaf_243_clk filters.res_lut\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_142_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17249_ _00319_ clknet_leaf_91_clk filters.sample_filtered\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09773__A1 _02131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11580__A1 _03673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08953_ _01411_ _01404_ _01417_ _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_110_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11707__I0 channels.atk_dec1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09525__A1 channels.sus_rel3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11637__I _03730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13321__A2 _04375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09525__B2 channels.pw2\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08884_ _01352_ _01353_ _01354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XPHY_EDGE_ROW_102_Left_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11332__A1 _03513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_2_clk_I clknet_5_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09505_ _01895_ _01896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12832__A1 _04831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_175_3627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_175_3638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09436_ _01782_ _00998_ _01827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_23_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15779__I _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09367_ filters.filt_3 _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_136_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_111_Left_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_164_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12596__B1 _04601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08681__I _01164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09298_ _01032_ _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_145_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14337__A1 _06211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16831__C _07710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11260_ _03202_ _03194_ _03201_ _03470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_105_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09764__A1 channels.atk_dec1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10211_ channels.pw1\[3\] _02430_ _02472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11191_ _03405_ _03389_ _03406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11571__A1 channels.freq3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10142_ _01085_ _02396_ _02393_ _02401_ _02402_ _02403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XTAP_TAPCELL_ROW_37_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10073_ _02319_ _02340_ _02343_ _00261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14950_ _01745_ channels.sample1\[0\] channels.sample2\[0\] _01759_ _06923_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_54_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16559__B _08339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13901_ _05900_ _05901_ _05902_ _05903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14881_ _06472_ _06820_ _06860_ _06861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15065__A2 _07033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13832_ _04397_ _04818_ _05835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_16620_ _08380_ _08384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13615__A3 _05220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16551_ _08314_ _08332_ _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_173_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13763_ _05671_ _05766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10975_ _03199_ _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15502_ filters.mode_vol\[7\] _01773_ _03214_ _03215_ _07444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_35_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12714_ _04366_ _04279_ _04720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_168_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16482_ _08237_ _08274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_168_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13694_ _04694_ _05075_ _05698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_5_0__f_clk clknet_3_0_0_clk clknet_5_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_38_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15433_ _07369_ _06910_ _07379_ _07381_ _06917_ _00583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_12645_ _04639_ _04640_ _04646_ _04650_ _04651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_150_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15364_ _07303_ _07304_ _07318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09452__B1 _01842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12576_ _04521_ _04527_ _04582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_81_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17103_ _00173_ clknet_leaf_110_clk channels.atk_dec1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__10062__A1 _02308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14328__A1 _05909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14315_ _06216_ _06228_ _06313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11527_ channels.pw1\[6\] _03650_ _03652_ _03655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15295_ _07203_ _07251_ _07254_ _07255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_17034_ _00104_ clknet_leaf_216_clk channels.lfsr\[1\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_150_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14246_ _06243_ _06244_ _06245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_22_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11458_ _03611_ _03603_ _01503_ _03604_ _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10409_ _02606_ _02609_ _02670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__12841__I _04220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14177_ _06066_ _06177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_11389_ channels.accum\[2\]\[9\] _03571_ _03572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_111_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13128_ _05115_ _05127_ _05133_ _05134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13059_ _04699_ _04221_ _04274_ _04511_ _05065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_178_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16253__A1 _07923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16818_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[1\] _00916_ _00918_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13067__A1 _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12288__I _04198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16749_ _00867_ _00868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_157_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08494__A1 filters.res_filt\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15820__C _07710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09221_ _01610_ _01659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_33_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09152_ _01594_ _01592_ _01598_ _01599_ _00080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_56_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_170_3535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_170_3546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10053__A1 channels.sus_rel3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09994__A1 channels.ctrl_reg3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09083_ _01323_ _01537_ _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_131_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09746__A1 _02112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10356__A2 _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_168_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09985_ channels.ctrl_reg3\[3\] _02276_ _02277_ _02281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_149_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08936_ _01400_ _01401_ _01402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__11305__A1 _01812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10108__A2 channels.ctrl_reg2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08867_ _01327_ _01329_ _01338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_157_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16244__A1 filters.sample_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13058__A1 _04699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08676__I _01159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13058__B2 _04697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08798_ channels.ctrl_reg3\[1\] channels.sync_outs\[1\] _01082_ _01271_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_54_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10760_ _02980_ _02981_ _03011_ _03015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_149_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09419_ _01811_ _01812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_164_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14558__A1 _05510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10292__A1 _02484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10691_ _02686_ _02923_ _02948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12430_ _04328_ _04363_ _04413_ _04436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_81_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_180_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10044__A1 channels.sus_rel3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16842__B _01753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09985__A1 channels.ctrl_reg3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11051__B _03273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12361_ _04366_ _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_106_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14100_ _06091_ _06099_ _06100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_95_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11312_ _03511_ _03508_ _03512_ _00331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_106_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15080_ _07044_ _07047_ _07048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_121_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12292_ _04292_ _04293_ _04296_ _04297_ _04298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_39_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14031_ _03397_ _04403_ _04881_ _06032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11243_ _03450_ _03444_ _03449_ _03454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_56_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12661__I _04632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14730__A1 _06722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10347__A2 _02607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11174_ _03386_ _03389_ _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_98_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10125_ _02385_ _02386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15982_ _07849_ _07862_ _07863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09970__I channels.pw3\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17721_ _00791_ clknet_leaf_61_clk tt_um_rejunity_sn76489.tone\[0\].gen.counter\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10056_ _02330_ _02331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14933_ _03730_ _04170_ _06907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17652_ _00722_ clknet_leaf_51_clk tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08586__I _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13049__A1 _04641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14864_ _06835_ _06843_ _06844_ _06845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16603_ _08374_ _08375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13815_ _05722_ _05723_ _05818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_58_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17583_ _00653_ clknet_leaf_33_clk spi_dac_i.spi_dat_buff_1\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14795_ _06779_ _06782_ _06783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_97_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16534_ _07355_ _08318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_35_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13746_ _05748_ _05749_ _05750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10958_ filters.filter_step\[0\] _03183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_161_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09673__B1 _01904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_223_clk_I clknet_5_20__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14549__A1 filters.band\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16465_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[7\] tt_um_rejunity_sn76489.tone\[2\].gen.counter\[6\]
+ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[5\] tt_um_rejunity_sn76489.tone\[2\].gen.counter\[4\]
+ _08259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_13677_ _05679_ _05638_ _05680_ _05681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11740__I _01150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10889_ _03127_ _03130_ _03132_ _03139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_14_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12628_ _04617_ _04634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15416_ _07364_ _07363_ _07365_ _07366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_16396_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[5\] _08201_ _08208_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12057__B _01032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15347_ _07290_ _07302_ _06979_ _00576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12559_ _03317_ _04506_ _04164_ _04565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_124_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_238_clk_I clknet_5_16__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15278_ _07202_ _07221_ _07238_ _07239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_124_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_112_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17017_ _00096_ clknet_leaf_229_clk channels.lfsr\[2\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14229_ _06219_ _06227_ _06228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14721__A1 filters.band\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_107_Right_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09770_ _02112_ _02125_ _02130_ _00171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08951__A2 _01415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_6_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15815__C _07269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08721_ _01174_ _01200_ _01204_ _01205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__09900__A1 channels.atk_dec2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08652_ channels.env_vol\[3\]\[7\] _01137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08496__I _01024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14788__A1 _06761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08583_ _01097_ _01098_ _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_77_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12746__I _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15122__I _06186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09204_ _01640_ _01641_ _01633_ _01642_ _01643_ _01644_ _01645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__15201__A2 _07122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16662__B _08339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10026__A1 _02289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09967__A1 _02250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09135_ _01583_ _01264_ _01095_ _01584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__14960__A1 filters.high\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09066_ _01519_ _01513_ _01521_ _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_128_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__16701__A2 _08437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13515__A2 _05520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12481__I _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11526__A1 _02324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11097__I _03316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09968_ channels.pw3\[10\] _02266_ _02262_ _02269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_51_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08919_ _01373_ _01371_ _01379_ _01386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09899_ _02150_ _02219_ _02221_ _00209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11930_ _04012_ _04013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16768__A2 net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10501__A2 _02754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11861_ _03748_ _03743_ _03950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13600_ _05471_ _05472_ _05605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10812_ _02955_ _02824_ _03066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14580_ _06425_ _06430_ _06575_ _06576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_0_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11792_ _03873_ _03874_ _03883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_135_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10265__A1 _01497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13531_ _05533_ _05535_ _05536_ _05537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_27_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10743_ _02992_ _02998_ _02999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_55_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16250_ _07923_ _08118_ _00663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13462_ _05314_ _05316_ _05467_ _05468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_11_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10674_ _02885_ _02931_ _02932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_40_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13203__A1 _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15201_ net56 _07122_ _07165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_35_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12413_ _04417_ _04418_ _04419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16181_ _08036_ _08052_ _08055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14871__I _05546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13393_ _05396_ _05397_ _05398_ _05399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_106_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15132_ _05404_ _07097_ _07098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_69_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12344_ _04252_ _04264_ _04350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_181_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15063_ _07007_ _07028_ _07031_ _07032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_121_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12275_ _04280_ _04281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11517__A1 channels.pw1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14014_ _04728_ _05347_ _06015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11226_ _03437_ _03434_ _03438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_71_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_243_clk clknet_5_5__leaf_clk clknet_leaf_243_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11157_ filters.high\[9\] _03373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__12317__I0 filters.cutoff_lut\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10108_ _01267_ channels.ctrl_reg2\[4\] _02369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15965_ _07813_ _07827_ _07846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11088_ _03297_ _03265_ _03266_ _03308_ _00311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_145_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17704_ _00774_ clknet_leaf_236_clk channels.lfsr\[0\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10039_ _02299_ _02310_ _02318_ _00252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_136_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14916_ filters.band\[30\] _03476_ _06892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15896_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[0\] _07766_ _07778_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__13690__A1 _05596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12493__A2 _04498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17635_ _00705_ clknet_5_23__leaf_clk channels.exp_counter\[0\]\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_69_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14847_ filters.band\[23\] _06820_ _06811_ _06830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_106_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_162_clk_I clknet_5_25__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17566_ _00636_ clknet_leaf_32_clk filters.low\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_86_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14778_ _06766_ _06767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_58_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16517_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[7\] _08270_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[7\]
+ _08304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_129_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_42_clk_I clknet_5_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13729_ _03350_ _04192_ _05732_ _05733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_17497_ _00567_ clknet_leaf_9_clk filters.high\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16448_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[2\] _08246_ _08098_ _08248_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_171_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16931__A2 _00923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10008__A1 channels.atk_dec3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_177_clk_I clknet_5_18__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09949__A1 _02215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13745__A2 _05657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14942__A1 _05534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16379_ _07809_ _08192_ _08193_ _08195_ _00715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_26_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_57_clk_I clknet_5_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_100_clk_I clknet_5_13__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_1308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09822_ _02137_ _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_165_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12308__I0 filters.cutoff_lut\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10192__C2 _01533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_115_clk_I clknet_5_26__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_182_3770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09753_ channels.ctrl_reg1\[5\] _02117_ _02113_ _02119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_182_3781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08704_ _01173_ _01188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09684_ filters.res_filt\[7\] _02007_ _02012_ channels.pw3\[7\] _02068_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_119_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08635_ _01128_ _00034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_167_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08566_ _01070_ _01082_ _01083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_37_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08497_ _01015_ _01026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_147_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_181_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14933__A1 _03730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09118_ _01562_ _01518_ _01568_ _01525_ _00077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_150_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10390_ _02612_ _02626_ _02650_ _02651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_32_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09049_ _01505_ _01506_ _01507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12060_ channels.env_counter\[0\]\[0\] _04108_ _04109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16438__A1 _08136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_225_clk clknet_5_20__leaf_clk clknet_leaf_225_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11011_ _03235_ _03236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_95_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11555__I _01812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12962_ _04486_ _04492_ _04968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_5_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15750_ _07661_ _07662_ _00619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12475__A2 _04480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11913_ _03906_ _03847_ _03911_ _03996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_14701_ filters.band\[11\] _05540_ _05541_ _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11683__B1 _03766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15681_ filters.sample_filtered\[14\] _07601_ _07610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12893_ _04823_ _04826_ _04899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_17420_ _00490_ clknet_leaf_137_clk channels.env_counter\[0\]\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11844_ _03934_ _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_14632_ _06623_ _06626_ _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09628__B1 _01964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13424__A1 _05289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10238__A1 _02484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17351_ _00421_ clknet_leaf_101_clk channels.freq3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12386__I _04258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14563_ _06542_ _06558_ _06559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11775_ channels.env_counter\[0\]\[4\] channels.env_counter\[1\]\[4\] channels.env_counter\[2\]\[4\]
+ channels.env_counter\[3\]\[4\] _03831_ _01167_ _03866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_32_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_101_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16302_ _08148_ _00685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13514_ _05515_ _05517_ _05519_ _05520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_10726_ _02980_ _02981_ _02982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_137_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17282_ _00352_ clknet_leaf_152_clk channels.accum\[2\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14494_ _06308_ _06388_ _06491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_81_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16913__A2 _03728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16233_ _08083_ _08104_ _08105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13445_ _05349_ _05352_ _05450_ _05451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__14924__A1 filters.band\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10657_ _02860_ _02861_ _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_181_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16164_ _07930_ _07850_ _07884_ _08039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_153_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13376_ _04911_ _05380_ _05381_ _05382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_10588_ _02802_ _02847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_50_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12327_ _03302_ _04332_ _04333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15115_ _07079_ _07081_ _07082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_16095_ _07954_ _07969_ _07972_ _07973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_107_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15046_ _07013_ _07014_ _07015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_103_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14152__A2 _05504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12258_ _04256_ _04260_ _04263_ _04264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_147_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_216_clk clknet_5_21__leaf_clk clknet_leaf_216_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_103_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11209_ filters.low\[12\] _03422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_12189_ _04194_ _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_143_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16997_ _00076_ clknet_leaf_189_clk channels.accum\[0\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_160_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15948_ _07810_ _07829_ _07830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13663__A1 _05584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12466__A2 _04468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15381__B _07333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15879_ _07760_ _07761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_121_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16601__A1 tt_um_rejunity_sn76489.chan\[1\].attenuation.in vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17618_ _00688_ clknet_leaf_139_clk channels.env_counter\[3\]\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13415__A1 _05417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10229__A1 _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12296__I _04207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13966__A2 _05967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17549_ _00619_ clknet_leaf_175_clk filters.low\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11977__A1 _04019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08842__A1 _01303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14766__I1 filters.band\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_119_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10952__A2 _01261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_160_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14143__A2 _06008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15340__A1 _07295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_207_clk clknet_5_20__leaf_clk clknet_leaf_207_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_61_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_180_3718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_3729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09805_ _02154_ _02155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__16840__A1 _06917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09736_ _02106_ _02107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_2_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09322__A2 _01734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09667_ _02048_ _02049_ _02050_ _02051_ _02052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_96_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08618_ channels.lfsr\[3\]\[13\] _01120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08684__I _01167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09598_ _01965_ _01973_ _01980_ _01985_ _01986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_167_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08549_ _01065_ clk_ctr\[1\] _01066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13957__A2 _05935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16834__C _04101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_1308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11560_ _03677_ _03669_ _03678_ _00413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09181__S1 _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10511_ _01668_ _02771_ _02772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14906__A1 _06456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13709__A2 _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11491_ _03513_ _03625_ _03630_ _00392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_52_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15310__I _06186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13230_ _03363_ _04271_ _04450_ _05236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_10442_ _02505_ _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_21_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12393__A1 _04200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13161_ _05066_ _05072_ _05167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10373_ _02519_ channels.env_vol\[3\]\[7\] _02633_ _02634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_60_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12112_ channels.accum\[3\]\[4\] _04138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15331__A1 _06919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13092_ _05058_ _05096_ _05097_ _05098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_12043_ _04068_ _04075_ _04097_ _00477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16920_ _00990_ _00854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09010__A1 _01468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13893__A1 _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12696__A2 _04480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16851_ _00937_ _00939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15802_ _07355_ _07700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_137_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16782_ _07909_ _00885_ _00891_ _00889_ _00815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12448__A2 _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13994_ _05988_ _05994_ _05995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_88_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10459__A1 _01164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15733_ _06078_ _07637_ _07650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12945_ _04935_ _04950_ _04951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_73_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15664_ _07587_ _07582_ _07593_ _07595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12876_ _04881_ _04882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_83_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17403_ _00473_ clknet_leaf_149_clk channels.env_counter\[1\]\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11408__B1 _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14615_ _03396_ _06508_ _06609_ _06610_ _00536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_11827_ _03831_ channels.env_counter\[3\]\[13\] _03918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15595_ _07530_ _07531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_56_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14070__A1 _06065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17334_ _00404_ clknet_leaf_89_clk channels.pw1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11758_ _03848_ _03849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14546_ _06435_ _06444_ _06541_ _06542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16347__B1 _01334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_153_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10631__A1 _02687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10709_ _02964_ _02965_ _02966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17265_ _00335_ clknet_leaf_70_clk tt_um_rejunity_sn76489.control_tone_freq\[1\]\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11689_ _01425_ _03780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_37_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14477_ _06472_ _06473_ _06379_ _06474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_126_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16216_ _08059_ _08068_ _08089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_153_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13428_ _05364_ _05373_ _05434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14373__A2 _06370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17196_ _00266_ clknet_leaf_78_clk clk_trg\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_16147_ _07994_ _08022_ _08023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13359_ _04420_ _05281_ _05365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10934__A2 _02932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16078_ _07761_ _07955_ _07762_ _07956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_80_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13333__B1 _04712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09001__A1 _01422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15029_ _03282_ _06968_ _06999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10242__S0 _01145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16822__A1 _01766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput2 addr[1] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_166_Left_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09521_ channels.ctrl_reg2\[1\] _01830_ _01834_ channels.freq3\[9\] _01911_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_36_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11742__S0 _03832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09452_ channels.atk_dec2\[0\] _01838_ _01842_ channels.pw3\[8\] _01843_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_91_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15389__A1 _07321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09383_ net6 _01782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13939__A2 _05796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10983__B _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_138_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10622__A1 channels.sample3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_173_3588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08910__S1 _01161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_173_3599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_175_Left_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_rebuffer31_I _04177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15561__A1 filters.sample_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14116__A2 _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09528__C1 _01871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08679__I _01162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11319__B _03517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09719_ _01751_ _02093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10991_ _03215_ _03216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_179_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12730_ _04733_ _04734_ _04735_ _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA_output22_I net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10449__I _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12661_ _04632_ _04667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_78_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09059__A1 _01422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11612_ _03689_ _03714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14400_ _03360_ _03221_ _06398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_61_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12592_ _04468_ _04597_ _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15380_ _07332_ _07333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_182_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_19__f_clk clknet_3_4_0_clk clknet_5_19__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_136_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11543_ _02298_ _03666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_14331_ _06326_ _06327_ _06328_ _06329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_52_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17050_ _00120_ clknet_leaf_230_clk channels.lfsr\[1\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14262_ _06008_ _06261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11474_ channels.accum\[1\]\[21\] _03590_ _03621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15552__A1 channels.sample2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16001_ _07788_ _07794_ _07881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_13213_ _04386_ _04180_ _04824_ _04791_ _05219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_10425_ _02562_ _02686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14193_ _06190_ _06191_ _06192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09973__I _02272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10916__A2 _03156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13144_ _04386_ _04791_ _05150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10356_ _02562_ _02502_ _02617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_59_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13075_ _04201_ _04758_ _05081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10912__I _02365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10287_ _02523_ _02546_ _02547_ _02548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__08589__I _01104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13866__A1 _05852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12026_ channels.env_counter\[1\]\[6\] _04085_ _04088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16903_ channels.exp_counter\[3\]\[0\] _00981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09534__A2 _01891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16804__A1 _01741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16834_ _08441_ _00925_ _03520_ _04101_ _00831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09922__B _02232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16765_ _01806_ _00869_ _00878_ _00811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13977_ _05903_ _05959_ _05978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_15716_ _07636_ _07637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12928_ _04877_ _04907_ _04933_ _04934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_76_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16696_ _08434_ _08436_ _01823_ _00791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_38_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15647_ _07577_ _07578_ _07579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12859_ _04200_ _04864_ _04865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_158_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15578_ _03326_ _07513_ _07514_ _06067_ _07515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_155_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17317_ _00387_ clknet_leaf_189_clk channels.accum\[1\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14529_ _06450_ _06468_ _06525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_154_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17248_ _00318_ clknet_leaf_85_clk filters.sample_filtered\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_116_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17179_ _00249_ clknet_leaf_76_clk channels.sus_rel3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_133_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15818__C _07710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09883__I _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10907__A2 _02973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15846__A2 _07728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08952_ _01416_ _01417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_122_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08883_ channels.freq2\[3\] _01275_ _01288_ channels.freq1\[3\] _01353_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_79_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11653__I _01319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09504_ _01836_ _01840_ _01895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_116_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_177_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12832__A2 _04833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09435_ _01785_ _01826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_66_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_3628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10269__I channels.ch3_env\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_175_3639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09366_ _01766_ _01767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_118_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12596__A1 _04297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12484__I _04489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09461__A1 filters.cutoff_lut\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09297_ _01722_ _01723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_145_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09461__B2 filters.cutoff_lut\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15534__A1 channels.sample3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15795__I _07683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_1193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10210_ _01582_ _02455_ channels.pw3\[3\] _02471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_162_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11190_ _03386_ _03405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_140_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10141_ channels.accum\[0\]\[22\] channels.accum\[1\]\[22\] channels.accum\[2\]\[22\]
+ channels.accum\[3\]\[22\] _01495_ _01496_ _02402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_30_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10072_ filters.cutoff_lut\[13\] _02341_ _02342_ _02343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_54_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12520__A1 _03317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13900_ _05813_ _05843_ _05902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14880_ _06762_ _06860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13831_ _05729_ _05734_ _05833_ _05834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13076__A2 _05080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17517__CLK clknet_5_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16550_ _08324_ _08331_ _08332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_58_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13762_ _05678_ _05763_ _05764_ _05765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_10974_ _03191_ _03194_ _03197_ _03198_ _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_69_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15501_ _03202_ _07443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_12713_ _04708_ _04717_ _04718_ _04719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16481_ _08265_ _08273_ _00739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13693_ _04230_ _05256_ _05697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15432_ _06934_ _07380_ _07381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12644_ _04618_ _04649_ _04650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15773__A1 filters.low\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12394__I _04184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12575_ _04577_ _04580_ _04581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_15363_ _07293_ _07294_ _07305_ _07317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_182_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09452__A1 channels.atk_dec2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09452__B2 channels.pw3\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17102_ _00172_ clknet_leaf_111_clk channels.atk_dec1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14314_ _06201_ _06215_ _06312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11526_ _02324_ _03649_ _03654_ _00403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__14328__A2 _05092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15525__A1 channels.sample2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15294_ _07238_ _07252_ _07253_ _07254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_40_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17033_ _00103_ clknet_leaf_216_clk channels.lfsr\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_78_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_150_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14245_ _04697_ _05687_ _06244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11457_ channels.accum\[1\]\[14\] _03611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09917__B _02232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_150_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10408_ _02667_ _02668_ _02669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_68_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14176_ _06168_ _06175_ _06176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_104_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11388_ _02974_ _03571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_111_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13127_ _05102_ _05114_ _05133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10339_ _02569_ _02600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09507__A2 _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13058_ _04699_ _04291_ _04511_ _04697_ _05064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09063__S0 _01139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_175_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17572__D _00642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12009_ _03737_ _04004_ _01032_ _04077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_79_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16817_ _01741_ _00915_ _00917_ _00910_ _00824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12569__I _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16748_ _08461_ _08442_ _08444_ _00867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_88_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_159_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_157_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16679_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[5\] _08244_ _08421_ _08422_
+ _08423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_159_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08494__A2 _01013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09220_ channels.lfsr\[2\]\[11\] _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_3_2_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09151_ _01589_ _01599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_170_3536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10589__B1 _02847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_170_3547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09082_ _01536_ _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_86_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_131_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11002__A1 filters.lp vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15819__A2 _07636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09984_ _02252_ _02275_ _02280_ _00235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_168_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08935_ channels.accum\[0\]\[7\] channels.accum\[1\]\[7\] channels.accum\[2\]\[7\]
+ channels.accum\[3\]\[7\] _01148_ _01163_ _01401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_08866_ _01299_ _01337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__16244__A2 _07722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08797_ _01264_ _01268_ _01269_ _01270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_28_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13058__A2 _04291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14694__I _06688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09682__A1 channels.ctrl_reg3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08485__A2 _01012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09682__B2 channels.ctrl_reg1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09418_ net14 _01811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10292__A2 _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10690_ _02945_ _02946_ _02947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__15755__A1 _07665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09349_ _01751_ _01752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13230__A2 _04271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12360_ _04323_ _04366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__15507__A1 _03194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11051__C _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11311_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[1\] _03509_ _03503_ _03512_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_106_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11792__A2 _03874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16414__I _08194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12291_ _04281_ _04297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_39_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14030_ _03382_ _04341_ _05107_ _06031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11242_ _03452_ _03453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_56_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14730__A2 _06712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09293__S0 _01604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11558__I _01817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11173_ filters.sample_filtered\[8\] _03366_ _03388_ _03389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_38_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10124_ _02383_ _02384_ _02385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_98_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15981_ _07861_ _07862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14494__A1 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17720_ _00790_ clknet_leaf_67_clk tt_um_rejunity_sn76489.tone\[0\].gen.counter\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10055_ _02289_ _01956_ _02330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_14932_ _06761_ _06905_ _06906_ _00557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17651_ _00721_ clknet_leaf_51_clk tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14863_ _06722_ _06839_ _06844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11293__I net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13049__A2 _05049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16602_ _01319_ _01587_ _08374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13814_ _05722_ _05723_ _05817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_17582_ _00652_ clknet_leaf_46_clk spi_dac_i.spi_dat_buff_1\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14794_ _06780_ _06781_ _06782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16533_ _08314_ _08317_ _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13745_ _05747_ _05657_ _05658_ _05749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__09673__A1 channels.ctrl_reg2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10957_ _03181_ _03182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09673__B2 _02056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16464_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[3\] tt_um_rejunity_sn76489.tone\[2\].gen.counter\[2\]
+ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[1\] tt_um_rejunity_sn76489.tone\[2\].gen.counter\[0\]
+ _08258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_128_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14549__A2 _04506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15746__A1 _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13676_ _05604_ _05637_ _05680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10888_ _02358_ _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_152_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15415_ filters.low\[23\] _06862_ _07365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_TAPCELL_ROW_152_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12627_ _04616_ _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16395_ _08206_ _08207_ _08200_ _00719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_26_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15346_ _06983_ _07301_ _07302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12558_ _04535_ _04537_ _04564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_108_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11509_ _03641_ _03643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_124_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12852__I _04739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15277_ _07236_ _07237_ _07220_ _07238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_12489_ _04466_ _04494_ _04495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_79_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17016_ _00095_ clknet_5_16__leaf_clk channels.lfsr\[2\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14228_ _06221_ _06226_ _06227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_1_clk_I clknet_5_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12732__A1 _04173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14159_ _06139_ _06158_ _06159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_42_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13683__I _05588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08539__I0 _01019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08720_ _01201_ _01202_ _01203_ _01188_ _01204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__16226__A2 _07924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08651_ _01136_ _00042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_90_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08582_ _01072_ _01098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_152_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_124_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09664__A1 channels.ch3_env\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_119_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09664__B2 channels.atk_dec1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11471__A1 _03612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09203_ _01606_ _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_91_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09416__A1 filters.bp vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13212__A2 _04444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09134_ _01582_ _01583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_72_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10026__A2 _01943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09967__A2 _02265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14960__A2 _06919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09065_ _01519_ _01513_ _01521_ _01522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_163_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_7_Left_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_115_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09275__S0 _01144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09967_ _02250_ _02265_ _02268_ _00230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_176_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_51_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08687__I _01170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08918_ _01384_ _01385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_99_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09898_ channels.atk_dec2\[4\] _02220_ _02217_ _02221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08849_ _01320_ _01321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10231__B _01469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15976__A1 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[0\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11860_ _03939_ _03948_ _03949_ _00442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10811_ _02994_ _02776_ _03065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11791_ _03878_ _03880_ _03882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_0_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12254__A3 _04259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13530_ filters.band\[0\] _03471_ _05536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10742_ _02993_ _02997_ _02998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_138_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13461_ _04269_ _04182_ _05465_ _05466_ _05467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_10673_ _02888_ _02930_ _02931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_clkbuf_5_18__f_clk_I clknet_3_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14400__A1 _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_173_Right_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_168_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_164_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15200_ _07163_ _07164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_153_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12412_ _04289_ _04304_ _04418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16180_ _07743_ _08053_ _08054_ _00657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_51_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13392_ _05394_ _05395_ _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_180_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15131_ _07053_ _05416_ _05421_ _07096_ _07097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_62_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12343_ _04252_ _04264_ _04349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12274_ _04279_ _04280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15062_ _07007_ _07028_ _07030_ _07031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09266__S0 _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12714__A1 _04366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11225_ _03431_ _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14013_ _05951_ _06012_ _06013_ _06014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_120_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_71_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11156_ filters.sample_filtered\[9\] _03372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12317__I1 filters.res_lut\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10107_ _01540_ _02361_ _02368_ _00270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15964_ _07841_ _07842_ _07844_ _07753_ _07845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_41_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11087_ _03305_ _03307_ _03308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_145_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17703_ _00773_ clknet_leaf_236_clk channels.lfsr\[0\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10038_ channels.sus_rel3\[3\] _02311_ _02312_ _02318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14915_ filters.low\[30\] _06891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_15895_ _07768_ _07777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09894__A1 channels.atk_dec2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13690__A2 _05597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17634_ _00704_ clknet_leaf_197_clk channels.exp_counter\[0\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14846_ _06804_ _06828_ _06829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_19_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17565_ _00635_ clknet_leaf_32_clk filters.low\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_86_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09646__A1 channels.freq1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14777_ _06765_ _06766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11751__I _01166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11989_ _04001_ _04059_ _04060_ _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__09646__B2 channels.pw3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16516_ _08265_ _08303_ _00744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13728_ _05731_ _05732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_14_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17496_ _00566_ clknet_leaf_9_clk filters.high\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09221__I _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16447_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[2\] _08246_ _08247_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_112_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13659_ _05570_ _05663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15195__A2 channels.sample1\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_140_Right_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16378_ _08194_ _08195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14942__A2 _06915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14283__B _06281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15329_ _07277_ _07280_ _07285_ _07286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_81_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17385__CLK clknet_5_31__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16695__A2 _08274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09891__I _01776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09821_ _02110_ _02163_ _02166_ _00186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_165_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10192__A1 _01541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11926__I _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_182_3760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09752_ _01801_ _02116_ _02118_ _00165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_182_3782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08703_ _01178_ _01187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09683_ filters.cutoff_lut\[16\] _01988_ _02009_ channels.ch3_env\[7\] _02067_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_94_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09885__A1 channels.atk_dec2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08634_ channels.lfsr\[3\]\[21\] _01128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09637__A1 channels.ctrl_reg2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08565_ _01081_ _01082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09637__B2 channels.atk_dec2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08496_ _01024_ _01025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_119_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_170_clk clknet_5_24__leaf_clk clknet_leaf_170_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_88_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_165_1225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14933__A2 _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12944__A1 _04938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12492__I _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09117_ _01300_ _01567_ _01568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09048_ channels.freq2\[15\] _01280_ _01293_ channels.freq1\[15\] _01506_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_130_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14697__A1 _06689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11010_ _03234_ _03235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12172__A2 _04177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_222_clk_I clknet_5_20__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09306__I _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09325__B1 _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12961_ _04486_ _04492_ _04967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_5_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09876__A1 channels.ctrl_reg2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14700_ _06692_ _06694_ _06695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11912_ _01584_ _03910_ _03995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15680_ _07600_ _07605_ _07609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_12892_ _04823_ _04826_ _04898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11683__B2 _03039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14631_ _06577_ _06624_ _06625_ _06626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11843_ _03856_ _03876_ _03896_ _03933_ _03934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__09628__A1 filters.lp vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09628__B2 channels.sus_rel1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13424__A2 _05377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17350_ _00420_ clknet_leaf_101_clk channels.freq3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10238__A2 _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14562_ _06549_ _06557_ _06558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_56_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11774_ _03836_ _03839_ _03864_ _03865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16301_ channels.env_counter\[3\]\[6\] _08148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_64_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13513_ _04850_ _05518_ _05519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17281_ _00351_ clknet_leaf_165_clk channels.accum\[2\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10725_ _02942_ _02970_ _02981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14493_ _06406_ _06409_ _06489_ _06490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_82_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_161_clk clknet_5_28__leaf_clk clknet_leaf_161_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_165_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16232_ _08082_ _08085_ _08104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_67_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13444_ _05446_ _05449_ _05353_ _05450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10656_ _02896_ _02913_ _02914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_152_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16163_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[3\] _07800_ _08038_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10915__I _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13375_ _04914_ _04932_ _05381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10587_ _02809_ _02814_ _02845_ _02846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_106_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15114_ _07052_ _07054_ _07080_ _07081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_23_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12326_ _04276_ _04332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_181_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16094_ _07929_ _07970_ _07971_ _07972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_133_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15045_ _06984_ _06992_ _07014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09925__B _02232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12257_ _04261_ _04262_ _04263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_147_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_147_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11208_ filters.sample_filtered\[12\] _03421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_12188_ _03189_ _03192_ _03195_ filters.high\[3\] _04194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_4
XPHY_EDGE_ROW_79_Left_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11139_ _03353_ _03356_ _03357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_16996_ _00075_ clknet_leaf_157_clk channels.accum\[0\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13112__A1 _04535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15947_ _07824_ _07828_ _07829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_92_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_160_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14860__A1 filters.band\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11674__A1 channels.sus_rel3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15878_ _07759_ _02347_ _07760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_25_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_121_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17617_ _00687_ clknet_leaf_150_clk channels.env_counter\[3\]\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_121_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10298__S _01144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14829_ filters.low\[22\] filters.band\[22\] _06073_ _06813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_118_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13415__A2 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11481__I _00389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10229__A2 _02473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17548_ _00618_ clknet_leaf_8_clk filters.low\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_88_Left_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_144_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_152_clk clknet_5_29__leaf_clk clknet_leaf_152_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_11_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16365__A1 channels.ch3_env\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17479_ _00549_ clknet_leaf_29_clk filters.band\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_157_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13718__A3 _05721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15837__B _07573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_97_Left_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09555__B1 _01943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_180_3719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11656__I _02721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09804_ _01805_ _02154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_157_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16668__B _01753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09735_ _01781_ _01941_ _02106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_2_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_179_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09666_ filters.hp _02014_ _01899_ channels.sus_rel1\[6\] _02051_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_59_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08617_ _01119_ _00025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09597_ channels.freq3\[11\] _01834_ _01862_ channels.pw2\[11\] _01984_ _01985_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__12209__A3 _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11417__A1 _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08548_ clk_trg\[1\] _01065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_46_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15798__I _07636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_181_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_143_clk clknet_5_27__leaf_clk clknet_leaf_143_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_119_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08479_ _01008_ _01009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_107_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10510_ _02386_ _02771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_174_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11490_ channels.freq1\[2\] _03626_ _03627_ _03630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_135_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10441_ _02699_ _02700_ _02701_ _02702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13590__A1 _04476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13160_ _05134_ _05165_ _05166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10372_ _01305_ _02632_ _02633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12111_ _04137_ _00505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_103_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13091_ _05086_ _05095_ _05097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_103_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09745__B _02113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_161_clk_I clknet_5_28__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12042_ channels.env_counter\[1\]\[13\] _04078_ _04097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09546__B1 _01862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13342__A1 _04265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09010__A2 _01470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_41_clk_I clknet_5_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16850_ _00937_ _00938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15095__A1 filters.high\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09036__I _01138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15801_ _06822_ _07697_ _07699_ _07269_ _00633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_102_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16781_ _02098_ _00886_ _00891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_176_clk_I clknet_5_18__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13993_ _05992_ _05993_ _05994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_99_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15732_ _05973_ _07632_ _07649_ _00614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_12944_ _04938_ _04949_ _04950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_clkbuf_leaf_56_clk_I clknet_5_8__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15663_ _07587_ _07582_ _07593_ _07594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_73_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12875_ _04880_ _04881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_158_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17402_ _00472_ clknet_leaf_150_clk channels.env_counter\[1\]\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_83_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14614_ _06186_ _06610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11826_ channels.env_counter\[2\]\[13\] _03917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_139_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15594_ filters.sample_buff\[6\] _07529_ _07530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_55_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17333_ _00403_ clknet_leaf_89_clk channels.pw1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_56_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14545_ _06438_ _06443_ _06541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_134_clk clknet_5_31__leaf_clk clknet_leaf_134_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11757_ _03846_ _03847_ _03848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_172_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15501__I _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17264_ _00334_ clknet_leaf_71_clk tt_um_rejunity_sn76489.control_tone_freq\[1\]\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10631__A2 _02840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10708_ _02962_ _02963_ _02965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_114_clk_I clknet_5_26__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14476_ _06254_ _06473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_114_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11688_ _03534_ _03778_ _03779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__12908__A1 _04831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16215_ _08078_ _08087_ _08088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_141_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13427_ _05364_ _05373_ _05433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17195_ _00265_ clknet_leaf_53_clk tt_um_rejunity_sn76489.noise\[0\].gen.signal_edge.previous_signal_state_0
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10639_ _02852_ _02853_ _02897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13581__A1 _04176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16146_ _07996_ _07999_ _08022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_148_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13358_ _05361_ _05362_ _05363_ _05364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_106_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_129_clk_I clknet_5_30__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12309_ _04314_ _04315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16077_ _07876_ _07955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13289_ _05267_ _05285_ _05294_ _05295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_114_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15028_ net38 _06970_ _06998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__10147__A1 channels.pw1\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10380__I _02522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10242__S1 _01159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput3 addr[2] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_16979_ _00058_ clknet_leaf_180_clk channels.accum\[0\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09520_ _01823_ _01910_ _00141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_36_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11647__A1 _02272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17573__CLK clknet_5_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11742__S1 _01171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09451_ _01841_ _01842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_148_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09382_ _01780_ _01781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_177_3670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13640__B _05643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_125_clk clknet_5_27__leaf_clk clknet_leaf_125_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__16338__A1 _03978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_138_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_138_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_3589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_1304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15561__A2 _07493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12375__A2 _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09528__C2 channels.freq3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11386__I _01240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09718_ _01742_ _02090_ _02092_ _00157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10990_ _03201_ _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_96_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09649_ _02028_ _02034_ _02035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_97_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12850__A3 _04192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12010__I _04077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12660_ _04594_ _04637_ _04628_ _04666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10861__A2 _02890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11611_ _03711_ _03713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_33_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_61_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_116_clk clknet_5_26__leaf_clk clknet_leaf_116_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12591_ _04596_ _04597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_38_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14330_ _04446_ _05367_ _06328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11542_ _03664_ _03658_ _03665_ _00408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_135_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14261_ _06144_ _06145_ _06260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_11473_ _03620_ _03615_ _01552_ _03616_ _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_16000_ _07748_ _07875_ _07877_ _07879_ _07880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_123_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13212_ _04485_ _04444_ _05218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10424_ _02684_ _02685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_151_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14192_ _06101_ _06161_ _06191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_104_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13143_ _04278_ _04780_ _05149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10355_ _02613_ _02614_ _02615_ _02616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_59_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09519__B1 net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08990__A1 channels.freq2\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08990__B2 channels.freq1\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13074_ _04401_ _05079_ _05080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_10286_ _02537_ _02545_ _02547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12025_ _04034_ _04084_ _04087_ _00469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16902_ _00980_ _00846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16833_ _08462_ _00925_ _00927_ _04101_ _00830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_16764_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[9\] _00873_ _00877_ _00878_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13976_ _05886_ _05898_ _05976_ _05977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15715_ _07635_ _07636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_12927_ _04911_ _04914_ _04932_ _04933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_16695_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[8\] _08274_ _08435_ _08436_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_29_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15646_ channels.sample1\[10\] _03428_ _07578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12858_ _04483_ _04864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_69_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11809_ _03898_ _03900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12054__A1 _03744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12855__I _04860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_107_clk clknet_5_15__leaf_clk clknet_leaf_107_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_7_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15577_ _01927_ _07488_ _07514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12789_ _03301_ _04314_ _04276_ _04795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__15791__A2 _07682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_155_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17316_ _00386_ clknet_leaf_156_clk channels.accum\[1\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_155_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14528_ _06453_ _06467_ _06524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09470__A2 _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17247_ _00317_ clknet_leaf_86_clk filters.sample_filtered\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_181_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14459_ filters.band\[29\] _06456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__16740__A1 _08453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_72_Right_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_153_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17178_ _00248_ clknet_leaf_122_clk channels.atk_dec3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_133_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16129_ _07981_ _08002_ _08005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_141_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12590__I _04529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08981__A1 _01442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08951_ _01414_ _01415_ _01416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08882_ channels.freq3\[3\] _01075_ _01352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_81_Right_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_5_25__f_clk clknet_3_6_0_clk clknet_5_25__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_179_3710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_16_Left_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_168_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09503_ channels.pw1\[8\] _01891_ _01893_ channels.freq2\[8\] _01894_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12293__A1 _04281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12832__A3 _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09434_ _01824_ _01825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_52_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_3629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09365_ _01765_ _01766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_23_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09296_ _01721_ _01722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_90_Right_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10359__A1 _01657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10140_ _02398_ _02399_ _02400_ _02401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_28_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10071_ _02334_ _02342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_54_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12520__A2 _04525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10531__A1 _02686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11844__I _03934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13830_ _05730_ _05733_ _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_98_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09314__I _01728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13761_ _05681_ _05740_ _05764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10973_ filters.band\[0\] _03198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_168_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15500_ _07436_ _06910_ _07441_ _07442_ _06917_ _00589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_12712_ _04701_ _04707_ _04718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16480_ _08262_ _08272_ _08273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_167_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13692_ _05595_ _05694_ _05695_ _05696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_35_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15222__A1 _01748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15431_ _07370_ _07371_ _07378_ _07380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_182_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12643_ _04594_ _04537_ _04648_ _04261_ _04649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__15773__A2 _07670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15362_ _07293_ _07305_ _07316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_12574_ _04565_ _04567_ _04579_ _04580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_109_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17101_ _00171_ clknet_leaf_112_clk channels.atk_dec1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14313_ _06309_ _06310_ _06311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11525_ channels.pw1\[5\] _03650_ _03652_ _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14890__I _06760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15293_ _07217_ _07237_ _07234_ _07253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_29_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17032_ _00102_ clknet_leaf_213_clk channels.lfsr\[1\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_78_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14244_ _04699_ _05505_ _06243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_150_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11456_ _03600_ _01487_ _03610_ _00377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_78_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_150_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10407_ _02653_ _02661_ _02663_ _02668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_14175_ _05877_ _06170_ _06174_ _06175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_11387_ _03568_ _03569_ _01420_ _03570_ _00348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__15289__A1 _05852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13126_ _05129_ _05130_ _05131_ _05132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_111_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10338_ _02598_ _02599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_42_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13057_ _04895_ _05061_ _05062_ _05063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_10269_ channels.ch3_env\[3\] _02530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09063__S1 _01480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12008_ _04075_ _04076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_84_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__16789__A1 _03499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16816_ _07801_ _00916_ _00917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16747_ _01806_ _08465_ _00866_ _00805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13959_ _05899_ _05960_ _05961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_177_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16678_ _08416_ _08420_ _08281_ _08422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15629_ filters.sample_buff\[8\] _07554_ _07562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_29_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13775__A1 _04764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09150_ _01595_ _01596_ _01593_ _01597_ _01140_ _01154_ _01598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_84_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_170_3537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_170_3548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09081_ _01526_ _01528_ _01534_ _01536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_182_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_131_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11929__I _04011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11002__A2 _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12750__A2 _04743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09983_ channels.ctrl_reg3\[2\] _02276_ _02277_ _02280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_168_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08934_ _01398_ _01399_ _01400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_42_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12502__A2 _04504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_24_Left_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08865_ channels.accum\[0\]\[2\] _01336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_97_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08796_ _01267_ channels.ctrl_reg3\[3\] channels.ctrl_reg1\[3\] _01252_ _01269_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_TAPCELL_ROW_28_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15452__A1 _07373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input14_I bus_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12266__A1 _03362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_154_Right_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09131__A1 _01270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09417_ _01807_ _01802_ _01810_ _00138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_109_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09348_ _01750_ _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_33_Left_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13230__A3 _04450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14924__B _06899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09279_ channels.lfsr\[1\]\[19\] _01708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_105_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15507__A2 _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11310_ _02184_ _03511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_22_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12290_ _04295_ _04296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_16_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11241_ filters.sample_filtered\[14\] _03452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_120_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09293__S1 _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09309__I _01730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08945__A1 _01400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11172_ _03387_ _03370_ _03388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_140_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_0__f_clk_I clknet_3_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10123_ channels.ctrl_reg2\[7\] _01273_ _01286_ channels.ctrl_reg1\[7\] _02384_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_15980_ _07855_ _07860_ _07861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09753__B _02113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_42_Left_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10054_ _02328_ _02320_ _02329_ _00256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14931_ filters.band\[31\] _04160_ _06775_ _06906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11701__C2 channels.atk_dec1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17650_ _00720_ clknet_leaf_51_clk tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14862_ _06840_ _06843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_16601_ tt_um_rejunity_sn76489.chan\[1\].attenuation.in _08370_ _08373_ _00759_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13813_ _05712_ _05814_ _05815_ _05816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_98_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17581_ _00651_ clknet_leaf_45_clk spi_dac_i.spi_dat_buff_1\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12257__A1 _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14793_ _06753_ _06757_ _06773_ _06781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_159_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_121_Right_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16532_ _08310_ _08316_ _08317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_98_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13744_ _05657_ _05658_ _05747_ _05748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10956_ filters.filter_step\[1\] _03181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_156_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09673__A2 _01830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16463_ _08241_ _08257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_112_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13675_ _05602_ _05679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_51_Left_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10887_ _03054_ _03136_ _03137_ _00281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_156_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15414_ _07363_ _06852_ _07364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_14_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12626_ _04619_ _04632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_182_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16394_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[5\] _08198_ _08207_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_152_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_152_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15345_ _07293_ _07300_ _07301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_124_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12557_ _04468_ _04562_ _04563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09928__B _02232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13509__A1 _04705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11508_ _03641_ _03642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15276_ _05751_ _07219_ _07237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_151_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12488_ _04475_ _04482_ net71 _04494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_110_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17015_ _00094_ clknet_leaf_238_clk channels.lfsr\[2\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_111_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14227_ _06222_ _06225_ _06226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_110_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11439_ _02364_ _03600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_106_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08936__A1 _01400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12732__A2 _04737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14158_ _06142_ _06157_ _06158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_1_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_60_Left_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_95_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13109_ _05102_ _05114_ _05115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_14089_ _06087_ _06088_ _06089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_95_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15682__A1 filters.sample_buff\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input6_I addr[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11484__I _03624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08650_ channels.env_vol\[3\]\[6\] _01136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_178_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08581_ _01096_ _01097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_17779_ _00849_ clknet_leaf_197_clk channels.exp_counter\[3\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_124_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09202_ _01604_ _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_147_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09133_ _01249_ _01582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_17_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09064_ _01520_ _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_114_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_90_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09966_ channels.pw3\[9\] _02266_ _02262_ _02268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_34_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15673__A1 filters.sample_buff\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08917_ _01377_ _01378_ _01384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_51_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09897_ _02209_ _02220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_96_clk clknet_5_13__leaf_clk clknet_leaf_96_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09352__A1 _01742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08848_ _01070_ _01319_ _01320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_169_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08779_ _01095_ _01252_ _01253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_58_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_108_Left_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_174_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09799__I _02149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13987__A1 _04630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10810_ _03028_ _02872_ _03064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_170_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11790_ _03878_ _03880_ _03881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_68_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10738__I _02638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10741_ _02995_ _02996_ _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_83_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13460_ _04805_ _05466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_137_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10672_ _02928_ _02929_ _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_11_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14400__A2 _03221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12411_ _04301_ _04416_ _04300_ _04417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_168_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13391_ _05388_ _05382_ _05384_ _05397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_62_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_20_clk clknet_5_3__leaf_clk clknet_leaf_20_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_63_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15130_ _05427_ _05428_ _07096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12342_ _04339_ _04347_ _04348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_63_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15061_ _07029_ _07030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_12273_ _04278_ _04279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09266__S1 _01680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14012_ _04694_ _05800_ _05256_ _05447_ _06013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__09039__I _01497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13911__A1 _04324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11224_ _03426_ _03429_ _03421_ _03436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_142_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_71_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09591__A1 _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11155_ _03358_ _03327_ _03328_ _03371_ _00315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_101_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10106_ channels.sync_outs\[0\] _01560_ _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15963_ _07761_ _07843_ _07844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11086_ filters.sample_filtered\[3\] _03291_ _03306_ _03307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_145_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_87_clk clknet_5_12__leaf_clk clknet_leaf_87_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_17702_ _00772_ clknet_leaf_236_clk channels.lfsr\[0\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_175_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10037_ _02316_ _02310_ _02317_ _00251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_145_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14914_ _06889_ _06890_ _00555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_15894_ _07773_ _07775_ _07776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_37_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17633_ _00703_ clknet_leaf_195_clk channels.exp_counter\[0\]\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_172_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14845_ _06825_ _06827_ _06828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_19_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17564_ _00634_ clknet_5_2__leaf_clk filters.low\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14776_ _06716_ _06765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_11988_ _03900_ _04058_ _04060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_86_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16515_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[6\] _08289_ _08300_ _08302_
+ _08303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_13727_ _04881_ _05731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_58_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10939_ channels.sample1\[5\] _03170_ _03171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17495_ _00565_ clknet_5_5__leaf_clk filters.high\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16446_ _04101_ _08245_ _08246_ _00731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_14_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13658_ _05577_ _05640_ _05661_ _05662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_45_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12609_ _04369_ _04615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_16377_ tt_um_rejunity_sn76489.noise\[0\].gen.restart_noise _01042_ _08194_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__11205__A2 _03403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13589_ _05515_ _05592_ _05593_ _05594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_82_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_11_clk clknet_5_7__leaf_clk clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_121_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15328_ _07278_ _07279_ _07285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15259_ _05751_ _07219_ _07220_ _07221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_41_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09820_ channels.freq2\[9\] _02164_ _02158_ _02166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_165_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15655__A1 filters.sample_buff\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14458__A2 _06261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09751_ channels.ctrl_reg1\[4\] _02117_ _02113_ _02118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_182_3761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_182_3772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_78_clk clknet_5_12__leaf_clk clknet_leaf_78_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_126_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08702_ _01185_ _01186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_94_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09682_ channels.ctrl_reg3\[7\] _01999_ _02004_ channels.ctrl_reg1\[7\] _02066_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_179_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08633_ _01127_ _00033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13969__A1 _03299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08564_ _01080_ _01081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_178_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08495_ _01010_ _01022_ _01023_ _01024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_0_147_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14394__A1 _06192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09116_ _01558_ _01566_ _01567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_44_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09270__B1 _01592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09047_ channels.freq3\[15\] _01080_ _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__10293__I _02553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14697__A2 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15646__A1 channels.sample1\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11380__B2 _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09949_ _02215_ _02247_ _02256_ _00224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_69_clk clknet_5_11__leaf_clk clknet_leaf_69_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_102_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09325__A1 _01689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13121__A2 _05121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12960_ _04505_ _04966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_5_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11911_ _03901_ _03922_ _03994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_169_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12891_ _04261_ _04896_ _04897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__11683__A2 _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14630_ _06578_ _06579_ _06625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_11842_ _03899_ _03901_ _03913_ _03932_ _03933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_135_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_0_clk_I clknet_5_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14561_ _06551_ _06556_ _06557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11773_ _03850_ _03845_ _03805_ _03864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11435__A2 _03593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16300_ _08147_ _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13512_ _04862_ _05518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_101_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17280_ _00350_ clknet_leaf_147_clk channels.accum\[2\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10724_ _02944_ _02969_ _02980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_64_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14492_ _06471_ _06488_ _06489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16231_ _08079_ _08086_ _08102_ _08103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13443_ _05448_ _05449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_81_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11818__S0 _01150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10655_ _02907_ _02912_ _02913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_64_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16162_ _07759_ _07982_ _07842_ _07877_ _08037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_3_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13374_ _04914_ _04932_ _05380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10586_ _02800_ _02808_ _02845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11299__I _02334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10946__A1 channels.sample1\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14137__A1 _06014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15113_ _03329_ _07051_ _07080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12325_ _04263_ _04329_ _04330_ _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_16093_ _07938_ _07942_ _07971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_11_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15044_ _06986_ _06991_ _07013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_12256_ filters.res_lut\[5\] _04168_ _04262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_147_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_147_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09564__A1 channels.pw3\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11207_ _03409_ _03392_ _03393_ _03420_ _00318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__09564__B2 channels.pw2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12187_ _03350_ _04187_ _04192_ _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_177_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11138_ filters.sample_filtered\[6\] _03337_ _03355_ _03356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_78_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_5_6__f_clk clknet_3_1_0_clk clknet_5_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_16995_ _00074_ clknet_leaf_161_clk channels.accum\[0\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13112__A2 _04896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09941__B _02243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15946_ _07825_ _07814_ _07827_ _07828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11069_ _03289_ _03290_ _03291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_0_clk clknet_5_4__leaf_clk clknet_leaf_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_160_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14860__A2 _04160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15877_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[3\] _07759_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_78_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17616_ _00686_ clknet_leaf_138_clk channels.env_counter\[3\]\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_121_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14828_ _06810_ _06812_ _00547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_121_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12218__A4 filters.high\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09175__S0 _01605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17547_ _00617_ clknet_leaf_242_clk filters.low\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14759_ _06732_ _06742_ _06749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_157_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17478_ _00548_ clknet_leaf_29_clk filters.band\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14376__A1 _06236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16429_ tt_um_rejunity_sn76489.control_noise\[0\]\[2\] tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[1\]
+ _08232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12593__I _04506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09555__A1 filters.cutoff_lut\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09555__B2 channels.sus_rel3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09803_ _02150_ _02151_ _02153_ _00181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_157_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09734_ _02104_ _02105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09858__A2 _01830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09665_ channels.freq1\[6\] _02011_ _02012_ channels.pw3\[6\] _02050_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11665__A2 _03531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08616_ channels.lfsr\[3\]\[12\] _01119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09596_ _01981_ _01982_ _01983_ _01984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_139_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09142__I _01590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08547_ clk_trg\[0\] _01063_ clk_ctr\[1\] _01064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_77_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_46_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08478_ filters.res_filt\[5\] _01005_ _01007_ _01008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_65_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10440_ _02697_ _02698_ _02701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_33_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09794__A1 channels.sus_rel1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13590__A2 _05077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10371_ channels.ch3_env\[7\] _02632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_61_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12110_ channels.accum\[3\]\[3\] _04137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13090_ _05086_ _05095_ _05096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_20_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09546__A1 channels.ctrl_reg3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12041_ _04064_ _04075_ _04096_ _00476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09546__B2 channels.pw2\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11353__A1 channels.ctrl_reg2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15619__A1 channels.sample1\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15763__B _07671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15095__A2 _07062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15800_ _06828_ _07698_ _07699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_176_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16780_ _07817_ _00885_ _00890_ _00889_ _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_13992_ _04498_ _05990_ _05993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_142_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12943_ _04940_ _04948_ _04949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_15731_ _05969_ _07633_ _07648_ _07649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15662_ filters.sample_buff\[11\] _07592_ _07593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12874_ _04879_ _04880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_87_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17401_ _00471_ clknet_leaf_137_clk channels.env_counter\[1\]\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_83_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11825_ channels.env_counter\[0\]\[13\] channels.env_counter\[1\]\[13\] _03886_ _03916_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14613_ _06403_ _06608_ _06609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_56_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11408__A2 _01245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15593_ _07527_ _07528_ _07529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_56_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17332_ _00402_ clknet_leaf_97_clk channels.pw1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_28_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14544_ _06538_ _06539_ _06540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11756_ _03805_ _03835_ _03847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__16347__A2 _01317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10707_ _02962_ _02963_ _02964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_17263_ _00333_ clknet_leaf_75_clk tt_um_rejunity_sn76489.control_tone_freq\[2\]\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14475_ _06380_ _06472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11687_ _03550_ _03755_ _03757_ _03777_ _03778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_153_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16214_ _08079_ _08086_ _08087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_126_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13426_ _05423_ _05431_ _05432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_4
X_17194_ _00264_ clknet_leaf_89_clk filters.cutoff_lut\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10638_ _02858_ _02863_ _02856_ _02896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__13030__A1 _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09785__A1 _01819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16145_ _07988_ _08018_ _08020_ _08021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_148_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13357_ _05247_ _05264_ _05363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_140_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10569_ _02792_ _02828_ _02829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__16613__I _08380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11592__A1 _03662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12308_ filters.cutoff_lut\[9\] filters.res_lut\[9\] _04217_ _04314_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_16076_ _07953_ _07948_ _07954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_84_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13288_ _05198_ _05266_ _05294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_114_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15027_ filters.low\[4\] _06993_ _06996_ _06997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_12239_ _04234_ _04239_ _04244_ _04245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__11344__A1 _03039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11895__A2 _03978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16283__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16978_ _00057_ clknet_leaf_186_clk channels.accum\[0\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_155_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_127_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput4 addr[3] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_56_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15929_ _07810_ _07811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12588__I _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16035__A1 _07880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09450_ _01839_ _01840_ _01841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_91_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09381_ _01779_ _01780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_176_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_177_3660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09897__I _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_177_3671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_221_clk_I clknet_5_21__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10083__A1 _01933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14349__A1 _06314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_138_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15010__A2 _06955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_160_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09776__A1 channels.atk_dec1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_236_clk_I clknet_5_16__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11583__A1 channels.freq3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16897__I0 _00966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09528__B2 channels.sus_rel2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09137__I _01585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16274__A1 filters.sample_buff\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15077__A2 channels.sample2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13627__A3 _05487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09717_ channels.pw1\[8\] _02091_ _02084_ _02092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12835__A1 _04732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09700__A1 channels.freq1\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08503__A2 _00129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09648_ _02030_ _02031_ _02032_ _02033_ _02034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_69_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09579_ filters.res_filt\[3\] _01844_ _01893_ channels.freq2\[11\] _01967_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_167_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11610_ _03711_ _03712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_26_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12590_ _04529_ _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_61_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10074__A1 filters.cutoff_lut\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11541_ channels.freq2\[2\] _03659_ _03660_ _03665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15001__A2 _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14260_ _06139_ _06158_ _06258_ _06259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_162_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11472_ channels.accum\[1\]\[20\] _03620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__15758__B _07648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13211_ _05211_ _05216_ _05217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09767__A1 _02110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10423_ _02599_ _02684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09756__B _02120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14191_ _06103_ _06160_ _06190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13142_ _04179_ _04800_ _05148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_10354_ _02593_ _02595_ _02615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_59_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_59_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09519__A1 _01873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13073_ _05078_ _05079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_76_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10285_ _02537_ _02545_ _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11326__A1 _01740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__16589__B _08339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12024_ channels.env_counter\[1\]\[5\] _04085_ _04087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16901_ _00971_ channels.exp_periods\[1\]\[4\] _00974_ _00980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_168_Right_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16832_ _03491_ _03496_ _00927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16763_ _02101_ _00877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13975_ _05889_ _05897_ _05976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_15714_ _03216_ _03730_ _03205_ _07635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12926_ _04922_ _04931_ _04932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_16694_ _08238_ _08429_ _08433_ _08435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_158_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14579__A1 _06420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15645_ channels.sample2\[10\] _03424_ _07576_ _03234_ _07577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_150_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12857_ _04400_ _04862_ _04863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_75_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11808_ _03857_ _03897_ _03898_ _03899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_173_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13251__A1 _04266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12788_ net63 _04195_ _04374_ _04794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_15576_ _07488_ _07513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10065__A1 filters.cutoff_lut\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_155_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17315_ _00385_ clknet_leaf_190_clk channels.accum\[1\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11739_ _03804_ _03829_ _03830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_16_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14527_ _06480_ _06521_ _06522_ _06523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_155_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17246_ _00316_ clknet_leaf_85_clk filters.sample_filtered\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13003__A1 _04996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14458_ _04600_ _06261_ _06455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13967__I filters.low\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09758__A1 channels.ctrl_reg1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13409_ _05409_ net66 _05414_ _05415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_17177_ _00247_ clknet_leaf_123_clk channels.atk_dec3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_142_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14389_ _06373_ _06386_ _06387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_141_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_133_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11565__A1 channels.freq3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_133_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16128_ _07743_ _08003_ _08004_ _00655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_51_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_161_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08981__A2 _01443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14503__A1 _03374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08950_ channels.accum\[0\]\[8\] channels.accum\[1\]\[8\] channels.accum\[2\]\[8\]
+ channels.accum\[3\]\[8\] _01148_ _01163_ _01415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_16059_ _07931_ _07936_ _07937_ _07938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_20_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08881_ _01350_ _01347_ _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_135_Right_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_179_3700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_179_3711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09502_ _01892_ _01893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_116_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12293__A2 _04291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16559__A2 _08282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09433_ _01001_ _01824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_63_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09364_ net10 _01765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_23_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13242__A1 _04255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13242__B2 _04471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09420__I _01812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_40_clk_I clknet_5_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09997__A1 _02242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09295_ _01282_ _01587_ _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_129_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_175_clk_I clknet_5_18__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_55_clk_I clknet_5_8__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11308__A1 _03499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10070_ _02330_ _02341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09516__A4 _01906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_102_Right_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_54_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_113_clk_I clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10531__A2 _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12021__I _04077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13760_ _05681_ _05740_ _05763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_10972_ _03196_ _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08488__A1 _01017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12711_ _04716_ _04717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13691_ _05596_ _05597_ _05695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_clkbuf_leaf_128_clk_I clknet_5_30__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15222__A2 channels.sample1\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15430_ _07370_ _07371_ _07378_ _07379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12642_ filters.res_lut\[0\] _04170_ _04648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10047__A1 channels.sus_rel3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15361_ _07313_ _07314_ _07315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12573_ _03302_ _04332_ _04578_ _04579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_17100_ _00170_ clknet_leaf_111_clk channels.atk_dec1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11524_ _02319_ _03649_ _03653_ _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14312_ _06230_ _06251_ _06310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15292_ _07217_ _07237_ _07234_ _07252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_151_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14243_ _06151_ _06152_ _06241_ _06242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_17031_ _00008_ clknet_leaf_177_clk filters.res_lut\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11455_ channels.accum\[1\]\[13\] _03605_ _03610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12691__I _04392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_150_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17563__CLK clknet_5_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_150_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_5_31__f_clk clknet_3_7_0_clk clknet_5_31__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10406_ _02603_ _02604_ _02667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14174_ _06173_ _06174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_150_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11386_ _01240_ _03570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_110_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15289__A2 _07233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13125_ _05101_ _05128_ _05131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10337_ _02592_ _02598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_111_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13056_ _04900_ _04905_ _05062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10268_ _01656_ _02529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_175_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09912__A1 channels.sus_rel2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12007_ _04074_ _04075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10199_ _01265_ _01263_ channels.pw2\[0\] _02460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_108_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16815_ _00914_ _00916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16746_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[9\] _00861_ _00863_ _00866_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09676__B1 _01964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13958_ _05903_ _05959_ _05960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_159_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_157_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12909_ _04855_ _04856_ _04915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13471__B _05476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16677_ _08416_ _08420_ _08421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_76_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13889_ _05793_ _05891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15628_ filters.sample_buff\[9\] _07448_ _07561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_158_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10038__A1 channels.sus_rel3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09979__A1 channels.ctrl_reg3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15559_ _07485_ _07497_ _07435_ _00593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_170_3538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09080_ _01526_ _01528_ _01534_ _01535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_142_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17229_ _00299_ clknet_leaf_174_clk channels.sample1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16801__I _00905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09982_ _02250_ _02275_ _02279_ _00234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_40_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08933_ channels.freq2\[7\] _01277_ _01289_ channels.freq1\[7\] _01399_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12502__A3 _04182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08864_ _01322_ _01333_ _01335_ _00056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08795_ _01267_ channels.ctrl_reg2\[3\] _01268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_28_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12266__A2 _04271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09416_ filters.bp _01803_ _01809_ _01810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09347_ _01062_ _01750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_168_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09278_ channels.lfsr\[0\]\[19\] _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_62_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14715__A1 _06298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_95_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11529__A1 channels.pw1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11240_ _03243_ _03446_ _03449_ _03245_ _03451_ _00320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10201__A1 channels.pw1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14940__B _06913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11171_ _03367_ _03387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_30_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10122_ channels.ctrl_reg3\[7\] _01073_ _02383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_73_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10053_ channels.sus_rel3\[7\] _02321_ _02322_ _02329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14930_ _06769_ _06903_ _06904_ _06905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__11701__B2 channels.atk_dec2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14861_ _06761_ _06841_ _06842_ _00550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_16600_ tt_um_rejunity_sn76489.chan\[1\].attenuation.in _08370_ _08318_ _08373_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13812_ _05713_ _05714_ _05815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_17580_ _00650_ clknet_leaf_44_clk spi_dac_i.spi_dat_buff_1\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14792_ _06756_ _06772_ _06765_ _06780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_16531_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[9\] _08315_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[9\]
+ _08316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09122__A2 _01560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11465__B1 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13743_ _05743_ _05746_ _05747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_10955_ filters.filter_step\[2\] _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_57_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16462_ _08136_ _07924_ _00737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_39_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13674_ _05666_ _05677_ _05678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10886_ channels.sample3\[10\] _03105_ _03137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_167_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15413_ filters.low\[24\] _07363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_12625_ _04630_ _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_14_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16393_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[4\] _08201_ _08206_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_152_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_152_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12556_ _04561_ _04562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15344_ _07277_ _07294_ _07299_ _07300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11507_ _03640_ _01885_ _03641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__13509__A2 _05074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12487_ _04484_ _04486_ _04492_ _04493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__14406__I _05543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15275_ _05752_ _07219_ _07236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17014_ _00093_ clknet_leaf_236_clk channels.lfsr\[2\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14226_ _06223_ _06224_ _06225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11438_ _03599_ _03591_ _01395_ _03592_ _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_105_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_246_clk clknet_5_0__leaf_clk clknet_leaf_246_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_106_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14157_ _06147_ _06156_ _06157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09944__B _02243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16621__I _08382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11369_ channels.accum\[2\]\[1\] _03559_ _03560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11940__A1 _04019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13108_ _05103_ _05109_ _05113_ _05114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_14088_ _05440_ _05980_ _05994_ _06088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_13039_ _05011_ _05012_ _05045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_28_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_128_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16631__A1 _01689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08580_ _01071_ _01096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17778_ _00848_ clknet_leaf_196_clk channels.exp_counter\[3\]\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16729_ tt_um_rejunity_sn76489.latch_control_reg\[2\] _08461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_53_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_141_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08872__A1 _01341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09201_ channels.lfsr\[3\]\[7\] _01642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_147_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09132_ _01082_ _01581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_173_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09063_ channels.accum\[0\]\[16\] channels.accum\[1\]\[16\] channels.accum\[2\]\[16\]
+ channels.accum\[3\]\[16\] _01139_ _01480_ _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_163_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12184__A1 _03239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09965_ _02245_ _02265_ _02267_ _00229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_34_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08916_ channels.accum\[0\]\[6\] _01383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09896_ _02209_ _02219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13684__A1 _04176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08847_ _01295_ _01319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_100_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13890__I _05891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08778_ _01251_ _01252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_170_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11998__A1 _04044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10740_ _02955_ _02623_ _02996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10671_ _02892_ _02927_ _02929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12410_ _04302_ _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_11_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13390_ _05394_ _05395_ _05396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_35_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12411__A2 _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16689__A1 _08333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12341_ _04346_ _04347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_90_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15060_ _06981_ _07029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_160_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12272_ _04277_ _04278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__15766__B _07671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_121_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14011_ _05512_ _05256_ _05448_ _05800_ _06012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_11223_ _03421_ _03392_ _03393_ _03435_ _00319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xclkbuf_leaf_228_clk clknet_5_17__leaf_clk clknet_leaf_228_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_121_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13911__A2 _05078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09764__B _02120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09040__A1 _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11154_ _03367_ _03370_ _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__15113__A1 _03329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_27__f_clk_I clknet_3_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10105_ _02366_ _02361_ _02367_ _00269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15962_ _07757_ _07754_ _07843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11085_ _03294_ _03278_ _03293_ _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17701_ _00771_ clknet_leaf_226_clk channels.lfsr\[0\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10036_ channels.sus_rel3\[2\] _02311_ _02312_ _02317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_145_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10489__A1 _02507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14913_ _06456_ _06869_ _06860_ _06890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_145_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15893_ _07774_ tt_um_rejunity_sn76489.chan\[1\].attenuation.in _07775_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_175_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11150__A2 _03366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17632_ _00702_ clknet_leaf_195_clk channels.exp_counter\[0\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14844_ _06815_ _06817_ _06826_ _06827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_19_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17563_ _00633_ clknet_5_0__leaf_clk filters.low\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14775_ _06759_ _06764_ _00542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11987_ _03900_ _04058_ _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11989__A1 _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16514_ _08296_ _08299_ _08301_ _08302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_169_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13726_ _03333_ _04522_ _05625_ _05730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_129_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17494_ _00564_ clknet_leaf_249_clk filters.high\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10938_ _01460_ _03170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08854__B2 channels.freq1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16445_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[1\] tt_um_rejunity_sn76489.noise\[0\].gen.counter\[0\]
+ _08240_ _08246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__14927__A1 _06720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13657_ _05579_ _05639_ _05661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10869_ _03109_ _03120_ _03121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_156_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15520__I _07446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12608_ _04613_ _04171_ _04614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16376_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[1\] _08191_ _08193_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_137_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13588_ _04848_ _04850_ _04945_ _05518_ _05593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_54_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15327_ filters.low\[17\] _06293_ _07283_ _07284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__08701__S1 _01172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12539_ _04536_ _04543_ _04544_ _04545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_170_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15352__A1 _07295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15258_ _05646_ _07190_ _07188_ _07220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_219_clk clknet_5_21__leaf_clk clknet_leaf_219_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_14209_ _05183_ _04819_ _06208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09674__B _01905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09031__A1 _01479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15189_ _07129_ _07153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_165_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11495__I _03624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09750_ _02106_ _02117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_182_3762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13666__A1 _04500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_182_3773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08701_ channels.exp_counter\[0\]\[2\] channels.exp_counter\[1\]\[2\] channels.exp_counter\[2\]\[2\]
+ channels.exp_counter\[3\]\[2\] _01175_ _01172_ _01185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_09681_ _02061_ _02062_ _02063_ _02064_ _02065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_08632_ channels.lfsr\[3\]\[20\] _01127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_146_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13418__A1 _05289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08563_ _01079_ _01080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14091__A1 _06004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08494_ filters.res_filt\[7\] _01013_ _01023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15591__A1 channels.sample2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09115_ _01562_ _01563_ _01564_ _01565_ _01140_ _01154_ _01566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_161_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09270__A1 _01577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_92_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09046_ _01494_ _01497_ _01504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09948_ channels.freq3\[11\] _02248_ _02255_ _02256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09325__A2 _01734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09879_ channels.ctrl_reg2\[7\] _02202_ _02206_ _02207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_172_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_5_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11763__S0 _03832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11910_ _03884_ _03885_ _03888_ _03993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_12890_ _04777_ _04896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__16071__A2 _07726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11841_ _03914_ _03907_ _03929_ _03931_ _03932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_68_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11772_ _03860_ _03862_ _03863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14560_ _06552_ _06555_ _06556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08836__A1 _01308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12632__A2 _04541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13511_ _04237_ _05516_ _05517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10723_ _02936_ _02977_ _02978_ _02979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__10643__A1 _02590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_64_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14491_ _06476_ _06487_ _06488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_55_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16230_ _08078_ _08087_ _08102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_82_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13442_ _05447_ _05448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10654_ _02908_ _02911_ _02912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_81_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11818__S1 _01166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16161_ _08013_ _08024_ _08035_ _08036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_13373_ _05098_ _05287_ _05379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_10585_ _02816_ _02826_ _02843_ _02844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15112_ _05416_ _07066_ _07078_ _07079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_12324_ _04256_ _04260_ _04330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16092_ _07938_ _07942_ _07970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_121_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12255_ _03288_ _04197_ _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_15043_ _06994_ _06995_ _07011_ _07012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_11206_ _03416_ _03419_ _03420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_147_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09564__A2 _01842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12186_ _04191_ _04192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_43_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11137_ _03354_ _03340_ _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16994_ _00073_ clknet_leaf_156_clk channels.accum\[0\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15945_ _07826_ tt_um_rejunity_sn76489.chan\[3\].attenuation.in _07827_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_11068_ filters.high\[3\] _03210_ _03290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_160_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_160_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10019_ channels.atk_dec3\[5\] _02302_ _02303_ _02305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15876_ _07757_ _07751_ _07758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_25_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17615_ _00685_ clknet_leaf_139_clk channels.env_counter\[3\]\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_149_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14827_ filters.band\[21\] _06785_ _06811_ _06812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_121_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14073__A1 _03299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_121_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09175__S1 _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17546_ _00616_ clknet_leaf_242_clk filters.low\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14758_ _05546_ _06748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13709_ _04452_ _04713_ _05713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09669__B _02036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17477_ _00547_ clknet_leaf_29_clk filters.band\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14689_ _06663_ _06682_ _06683_ _06684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_144_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16428_ _08230_ _08231_ _08195_ _00728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_132_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14376__A2 _06249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12387__A1 _04392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16359_ channels.ch3_env\[2\] _08179_ _08182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10937__A2 _02973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09802_ channels.sus_rel1\[4\] _02152_ _02146_ _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_157_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09733_ _01739_ _02104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_66_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_2_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_2_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09664_ channels.ch3_env\[6\] _02009_ _01948_ channels.atk_dec1\[6\] _02049_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12862__A2 _04846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08615_ _01118_ _00024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_96_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09595_ filters.cutoff_lut\[12\] _01956_ _01954_ channels.freq1\[3\] _01983_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_49_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14064__A1 _06062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08546_ clk_ctr\[0\] _01063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_38_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12614__A2 _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11673__I0 _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08477_ _01006_ _01005_ _01007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_175_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15564__A1 channels.sample2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_149_Right_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10370_ _02598_ _02630_ _02576_ _02631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__14119__A2 _04927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09029_ _01422_ _01487_ _01488_ _00068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12040_ channels.env_counter\[1\]\[12\] _04078_ _04096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11353__A2 _01282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13991_ _05942_ _05944_ _05991_ _05992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_176_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15730_ _07355_ _07648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_172_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12942_ _04941_ _04944_ _04947_ _04948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_88_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12853__A2 _04858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_66_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15661_ _07590_ _07591_ _07592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14055__A1 _06024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12873_ filters.cutoff_lut\[15\] _04441_ _04879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_17400_ _00470_ clknet_leaf_139_clk channels.env_counter\[1\]\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_83_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14612_ _06602_ _06607_ _06608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_157_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11824_ _03890_ _03868_ _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_83_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13802__A1 _04728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15592_ channels.sample1\[6\] _03401_ _07528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17331_ _00401_ clknet_leaf_86_clk channels.pw1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14543_ _06458_ _06466_ _06539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11755_ _03845_ _03835_ _03846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17262_ _00332_ clknet_leaf_75_clk tt_um_rejunity_sn76489.control_tone_freq\[2\]\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15555__A1 filters.sample_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10706_ _02676_ _02824_ _02963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14474_ _06412_ _06470_ _06471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_113_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11686_ _03761_ _03764_ _03773_ _03776_ _03777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_181_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16213_ _08082_ _08085_ _08086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_36_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13425_ _05424_ _05425_ _05426_ _05429_ _05430_ _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_180_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17193_ _00263_ clknet_leaf_89_clk filters.cutoff_lut\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_23_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10637_ _02893_ _02875_ _02894_ _02895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_180_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10919__A2 _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16144_ _07988_ _08019_ _08020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_116_Right_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10568_ _02794_ _02827_ _02828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_24_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13356_ _05247_ _05264_ _05362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_3_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08840__C _01159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12307_ _04312_ _04313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_51_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16075_ _07943_ _07946_ _07953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13287_ _05274_ _05290_ _05292_ _05293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10499_ _02758_ _02759_ _02760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15026_ _06994_ _06995_ _06996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_114_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12238_ _03273_ _04243_ _04231_ _04244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XPHY_EDGE_ROW_126_Left_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__16807__A1 _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12169_ _04174_ _04175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16977_ _00056_ clknet_leaf_182_clk channels.accum\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14294__A1 _03347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput5 addr[4] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_36_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15928_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\] _07809_ _07810_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_36_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09170__B1 _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15859_ _07741_ _07742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_149_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09380_ _01003_ _01779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_135_Left_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_177_3661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_177_3672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17529_ _00599_ clknet_leaf_82_clk filters.sample_buff\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09473__A1 _01852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11280__A1 _02314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_138_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15546__A1 filters.sample_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14349__A2 _06346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11948__I _04006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10852__I _02974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_144_Left_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_125_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09418__I net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_168_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_7_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10138__A3 channels.pw3\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16274__A2 _07742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14285__A1 _03345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09716_ _02089_ _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11099__A1 filters.high\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09647_ filters.bp _02014_ _01964_ channels.sus_rel1\[5\] _02033_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_179_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_153_Left_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14037__A1 _05469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09578_ _01837_ _01966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_136_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12599__A1 _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08529_ _01050_ _00130_ _01052_ _01053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_182_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16915__S _00987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11540_ _01765_ _03664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_136_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15537__A1 channels.sample1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11471_ _03612_ _01545_ _03619_ _00383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_80_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10422_ _02669_ _02674_ _02681_ _02682_ _02683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_13210_ _05212_ _05215_ _05216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_150_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14190_ _06089_ _06100_ _06188_ _06189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XPHY_EDGE_ROW_162_Left_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_122_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12771__A1 filters.cutoff_lut\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10353_ _02593_ _02595_ _02614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13141_ _05143_ _05144_ _05146_ _05147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XTAP_TAPCELL_ROW_59_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09519__A2 _01889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13072_ _05077_ _05078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11079__B _03299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10284_ _02524_ _02543_ _02544_ _02545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_108_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12023_ _04029_ _04084_ _04086_ _00468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16900_ _00979_ _00845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16831_ _08443_ _00925_ _00926_ _07710_ _00829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_75_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16762_ _01800_ _00869_ _00876_ _00810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13974_ _05543_ _05975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_171_Left_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09152__B1 _01598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15713_ _05539_ _07632_ _07634_ _00610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_12925_ _04925_ _04928_ _04930_ _04931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_87_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16693_ _08280_ _08429_ _08433_ _08434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__09998__I _01779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10002__I _02174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15644_ _03409_ _07563_ _07575_ _03424_ _07576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_12856_ _04861_ _04862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_68_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11807_ channels.env_counter\[0\]\[11\] channels.env_counter\[1\]\[11\] channels.env_counter\[2\]\[11\]
+ channels.env_counter\[3\]\[11\] _01150_ _01165_ _03898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_15575_ filters.sample_buff\[4\] _07504_ _07512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_90_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12787_ _03315_ _04323_ net59 _04793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_83_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17314_ _00384_ clknet_leaf_157_clk channels.accum\[1\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14526_ _06484_ _06254_ _06483_ _06522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11738_ _03816_ _03827_ _03828_ _03829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_155_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_155_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17245_ _00315_ clknet_leaf_90_clk filters.sample_filtered\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14457_ filters.band\[28\] _05446_ _06454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_180_Left_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_172_3580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11669_ _03540_ _03759_ _03760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_116_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13408_ net61 _05412_ _05414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_98_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17176_ _00246_ clknet_leaf_123_clk channels.atk_dec3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_142_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14388_ _06376_ _06385_ _06386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14751__A2 _06703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12762__A1 _04714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16127_ spi_dac_i.spi_dat_buff_1\[4\] _07867_ _07921_ spi_dac_i.spi_dat_buff_1\[5\]
+ _03734_ _08004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_133_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13339_ _05342_ _05343_ _05344_ _05345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_84_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09238__I _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16058_ _07896_ _07902_ _07898_ _07937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14503__A2 _06177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15009_ _06956_ _06977_ _06979_ _00561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08880_ _01341_ _01342_ _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14267__A1 _05440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_179_3701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_179_3712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09501_ _01826_ _01836_ _01828_ _01892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_78_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09694__A1 _01742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13490__A2 _05345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09432_ _01822_ _01823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_52_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09363_ _01757_ _01743_ _01764_ _00126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_23_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13242__A2 _04864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09294_ _01716_ _01591_ _01720_ _01589_ _00101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_129_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_10 _01590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16534__I _07355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15578__C _06067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08957__B1 _01420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17365__CLK clknet_5_25__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11627__B _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16709__I _08445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09685__A1 channels.pw1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10971_ _03195_ _03196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_168_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12710_ _04709_ _04714_ _04715_ _04716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_167_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11492__A1 channels.freq1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15758__A1 _03422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output20_I net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13690_ _05596_ _05597_ _05694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_97_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12641_ _04639_ _04640_ _04646_ _04647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_167_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14430__A1 _04805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15360_ filters.low\[20\] _06599_ _07314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_148_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12572_ _04525_ _04578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_81_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15769__B _07671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14311_ _06197_ _06229_ _06309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11523_ channels.pw1\[4\] _03650_ _03652_ _03653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_124_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15291_ _07235_ _07221_ _07251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17030_ _00007_ clknet_5_18__leaf_clk filters.res_lut\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14242_ _04575_ _05774_ _06153_ _06241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_80_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11454_ _03609_ _03603_ _01475_ _03604_ _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_68_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_78_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_150_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_150_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10405_ _02653_ _02664_ _02665_ _02666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14173_ _06063_ _06171_ _06172_ _06173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_11385_ _01089_ _03569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_110_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_132_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13124_ _05060_ _05063_ _05083_ _05130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_10336_ _02585_ _02596_ _02597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_111_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13055_ _04900_ _04905_ _05061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10267_ _02527_ _02528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_12006_ _02363_ _04005_ _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_clkbuf_leaf_220_clk_I clknet_5_21__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15009__B _06979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10198_ _01498_ _02458_ _02459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16814_ _00914_ _00915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_17_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16745_ _01800_ _08465_ _00865_ _00804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_89_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13957_ _05905_ _05935_ _05958_ _05959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__09676__A1 channels.sus_rel3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09676__B2 channels.sus_rel1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12908_ _04831_ _04912_ _04913_ _04914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_clkbuf_leaf_235_clk_I clknet_5_16__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16676_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[5\] _08399_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[5\]
+ _08420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15749__A1 _03374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_157_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13888_ _04561_ _05883_ _05890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_158_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15627_ _07498_ _07560_ _00598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_174_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09428__A1 filters.mode_vol\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12839_ _04792_ _04796_ _04845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_174_3620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15558_ _07486_ _07495_ _07496_ _07497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_17_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14509_ _06502_ _06505_ _06506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_86_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_170_3539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15489_ net67 _07432_ _06952_ _07433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_182_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17228_ _00298_ clknet_leaf_176_clk channels.sample1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_142_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09287__S0 _01145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12735__A1 _04184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17159_ _00229_ clknet_leaf_121_clk channels.pw3\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_130_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09600__A1 _01933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10210__A2 _02455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09981_ channels.ctrl_reg3\[1\] _02276_ _02277_ _02279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_149_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08932_ channels.freq3\[7\] _01397_ _01398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08863_ channels.accum\[0\]\[1\] _01334_ _01335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_157_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08794_ _01266_ _01267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_58_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09667__A1 _02048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09431__I _01821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09415_ _01808_ _01809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11182__B _03396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13215__A2 _05220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09346_ _01013_ _01749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_118_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09277_ channels.lfsr\[2\]\[20\] _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11170_ filters.sample_filtered\[9\] _03385_ _03386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_56_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10121_ _02381_ _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_73_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14512__I _05544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10052_ _01818_ _02328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_14860_ filters.band\[24\] _04160_ _06775_ _06842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13811_ _05713_ _05714_ _05814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_138_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14791_ _06777_ _06778_ _06779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__09658__B2 channels.freq2\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16530_ _08242_ _08270_ _08315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13742_ _05555_ _05744_ _05745_ _05746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_39_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10954_ filters.sample_filtered\[0\] _03179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_39_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09341__I filters.filt_1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16461_ _08136_ _08256_ _00736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_97_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13673_ _05669_ _05676_ _05677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10885_ _03125_ _03135_ _03136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
Xclkbuf_leaf_191_clk clknet_5_22__leaf_clk clknet_leaf_191_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__14403__A1 _06298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15412_ _07340_ _07358_ _07359_ _07321_ _07361_ _07362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_12624_ _04629_ _04630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_66_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16392_ _08204_ _08205_ _08200_ _00718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_155_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15499__B _06913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12965__A1 _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15343_ _07297_ _07298_ _07299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_170_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12555_ _04500_ _04561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_93_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09830__A1 _02150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11506_ _01779_ _03640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_136_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15274_ _07225_ _07234_ _07235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_12486_ _04487_ _04491_ _04492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17013_ _00092_ clknet_leaf_238_clk channels.lfsr\[2\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14225_ _04893_ _05447_ _06224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_130_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11437_ channels.accum\[1\]\[6\] _03599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_111_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14156_ _06150_ _06155_ _06156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_81_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11368_ _02974_ _03559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_120_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13107_ _05110_ _05111_ _05112_ _05113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_21_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10319_ _01306_ channels.env_vol\[3\]\[5\] _02579_ _02580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_42_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14087_ _04645_ _06086_ _05992_ _06087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11299_ _02334_ _03503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_167_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13038_ _04952_ _04991_ _05044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_119_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_128_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_174_clk_I clknet_5_24__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14989_ _06943_ _06960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_17777_ _00847_ clknet_leaf_195_clk channels.exp_counter\[3\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11456__A1 _03600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16728_ _01806_ _08447_ _08460_ _00799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_54_clk_I clknet_5_10__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_141_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16659_ _08394_ _08404_ _08405_ _08406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_48_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_182_clk clknet_5_19__leaf_clk clknet_leaf_182_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_151_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08872__A2 _01342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09200_ channels.lfsr\[1\]\[7\] _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_53_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_189_clk_I clknet_5_22__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09131_ _01270_ _01579_ _01580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_69_clk_I clknet_5_11__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09821__A1 _02110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09062_ _01505_ _01506_ _01510_ _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__16698__A2 _08437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_112_clk_I clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12708__A1 _04186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11392__B1 _01448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_90_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_127_clk_I clknet_5_27__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09964_ channels.pw3\[8\] _02266_ _02262_ _02267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09426__I _01817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13133__A1 _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08915_ _01322_ _01381_ _01382_ _00060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09895_ _02215_ _02210_ _02218_ _00208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_51_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14881__A1 _06472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08846_ _01260_ _01262_ _01316_ _01318_ _00055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11695__B2 channels.atk_dec2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08777_ _01249_ _01250_ _01251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_79_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14633__A1 _04318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_173_clk clknet_5_24__leaf_clk clknet_leaf_173_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_178_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_49_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08863__A2 _01334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10100__I _01282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10670_ _02892_ _02927_ _02928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_168_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12947__A1 _04475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09329_ _01698_ _01736_ _01737_ _01574_ _00119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_11_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_168_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12340_ _04345_ _04340_ _04346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_168_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12271_ _03301_ _04276_ _04277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_65_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14010_ _06006_ _06010_ _06011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__13372__A1 _05289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11222_ _03431_ _03434_ _03435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_120_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10186__A1 _01533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11153_ filters.sample_filtered\[7\] _03352_ _03369_ _03370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09336__I net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10104_ channels.sync_outs\[1\] _01230_ _02367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15961_ _07747_ _07752_ _07842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11084_ filters.sample_filtered\[4\] _03304_ _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09879__A1 channels.ctrl_reg2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10035_ _02187_ _02316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_17700_ _00770_ clknet_leaf_226_clk channels.lfsr\[0\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14912_ _06851_ _06888_ _06889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_175_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10489__A2 _02512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15892_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[1\] _07774_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_145_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08551__A1 clk_trg\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08551__B2 clk_trg\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12697__I _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17631_ _00701_ clknet_leaf_204_clk channels.env_vol\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14843_ _06720_ _06813_ _06826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__14624__A1 _06520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17562_ _00632_ clknet_leaf_30_clk filters.low\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11438__B2 _03592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14774_ filters.band\[16\] _06761_ _06763_ _06764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11986_ _04053_ _04054_ _04058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_58_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16513_ _08257_ _08301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_123_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_86_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13725_ _04274_ _04819_ _05729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17493_ _00563_ clknet_leaf_6_clk filters.high\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10937_ _03168_ _02973_ _03169_ _00299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_164_clk clknet_5_28__leaf_clk clknet_leaf_164_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_128_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16444_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[0\] _08244_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[1\]
+ _08245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_39_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13656_ _05565_ _05576_ _05659_ _05660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_67_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10868_ _03116_ _03119_ _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_6_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12607_ _03256_ _04566_ _04613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_16375_ _08191_ _08192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_155_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10945__I _01320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09803__A1 _02150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13587_ _04238_ _04945_ _05518_ _04847_ _05592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10799_ _02882_ _03052_ _03053_ _00277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_30_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_136_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15326_ filters.low\[16\] _06287_ _07283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_170_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12538_ _04540_ _04542_ _04544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_83_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16632__I _08380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15257_ _07217_ _07218_ _07219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_12469_ _04387_ _04472_ _04474_ _04475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_83_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14208_ _06205_ _06206_ _06207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__12166__A2 _04171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15188_ _07125_ _07150_ _07151_ _07152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09031__A2 _01482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14139_ _06137_ _06138_ _06139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_165_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14863__A1 _06722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_182_3774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08700_ _01169_ _01183_ _01184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_182_3785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11677__A1 _01168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09680_ channels.atk_dec2\[7\] _01838_ _01937_ channels.freq3\[7\] _02064_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08631_ _01126_ _00032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13418__A2 _05377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14615__A1 _03396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_179_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08562_ _01078_ _01079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_178_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09098__A2 _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16368__A1 _03974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08493_ net15 _01011_ _01022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10101__A1 _01070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_155_clk clknet_5_29__leaf_clk clknet_leaf_155_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_77_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15711__I _07630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12229__I0 filters.cutoff_lut\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15040__A1 _05969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15591__A2 _06397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09114_ channels.accum\[3\]\[22\] _01565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11601__A1 _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_92_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09045_ _01489_ _01409_ _01503_ _01421_ _00069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_103_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09947_ _02254_ _02255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_110_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11668__A1 channels.sus_rel3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09878_ _02175_ _02206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11668__B2 channels.sus_rel2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11763__S1 _03842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08829_ channels.freq2\[0\] _01274_ _01287_ channels.freq1\[0\] _01302_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__14606__A1 _06599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11840_ _03930_ _03931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12310__I _04315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11771_ _03861_ _03862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_146_clk clknet_5_28__leaf_clk clknet_leaf_146_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__16359__A1 channels.ch3_env\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13510_ _04740_ _05516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10722_ _02937_ _02971_ _02978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14490_ _06479_ _06486_ _06487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_101_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13441_ _05260_ _05447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10653_ _02909_ _02910_ _02911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_152_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15582__A2 _07518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16160_ _08034_ _08035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_51_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13372_ _05289_ _05377_ _05378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_181_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10584_ _02797_ _02815_ _02843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_106_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15111_ filters.low\[7\] _07077_ _07078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_134_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12323_ _04256_ _04260_ _04329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16091_ _07956_ _07958_ _07968_ _07969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_23_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_39_Left_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__15334__A2 _06955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_181_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09549__B1 _01937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15042_ _05014_ _05046_ _04993_ _07011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_107_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12254_ _03272_ _04243_ _04259_ _04260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_146_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11205_ filters.sample_filtered\[10\] _03403_ _03418_ _03419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_103_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_147_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12185_ _04190_ _04191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15098__A1 _05417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11136_ _03338_ _03354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_78_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16993_ _00072_ clknet_leaf_192_clk channels.accum\[0\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15944_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[0\] _07826_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_11067_ _03282_ _03188_ _03288_ _03206_ _03289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_125_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_160_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10018_ _02234_ _02301_ _02304_ _00245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_160_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15875_ _07756_ _07757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_48_Left_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_17614_ _00684_ clknet_leaf_139_clk channels.env_counter\[3\]\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14826_ _06762_ _06811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_121_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14073__A2 _06073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15270__A1 _07227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17545_ _00615_ clknet_leaf_242_clk filters.low\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14757_ _06739_ _06508_ _06747_ _06610_ _00541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xclkbuf_leaf_137_clk clknet_5_31__leaf_clk clknet_leaf_137_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_153_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11969_ _04001_ _04044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__16627__I _08382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13708_ _04325_ _04924_ _05712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17476_ _00546_ clknet_leaf_245_clk filters.band\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14688_ _06543_ _06548_ _06546_ _06683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_157_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16427_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[14\] _08197_ _08231_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13639_ _05549_ _05550_ _05643_ _05644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_0_128_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13584__A1 _04400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16358_ _03948_ _08177_ _08181_ _00708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_57_Left_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15309_ _07265_ _07266_ _07267_ _07268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_171_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16289_ channels.env_counter\[3\]\[0\] _08142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_180_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13336__A1 _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15089__A1 _03310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09801_ _02141_ _02152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09732_ _02097_ _02090_ _02099_ _02103_ _00160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__13654__C _05643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09663_ filters.res_filt\[6\] _02007_ _01939_ channels.sample3\[10\] _02048_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_2_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10322__A1 _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08614_ channels.lfsr\[3\]\[11\] _01118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_179_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09594_ channels.atk_dec3\[3\] _01867_ _01895_ channels.pw3\[3\] _01982_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08545_ net17 _01062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xclkbuf_leaf_128_clk clknet_5_30__leaf_clk clknet_leaf_128_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__13811__A2 _05714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08476_ net13 _01006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_119_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15564__A2 _03377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09028_ channels.accum\[0\]\[13\] _01461_ _01488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10561__A1 _01689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14827__A1 filters.band\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13990_ _04616_ _05990_ _05945_ _05991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_142_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12941_ _04416_ _04946_ _04947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15660_ channels.sample1\[11\] _03428_ _07591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12872_ _04821_ _04827_ _04878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_103_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14055__A2 _06055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14611_ _06298_ _06603_ _06606_ _06607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_11823_ _03905_ _03914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_83_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_119_clk clknet_5_26__leaf_clk clknet_leaf_119_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_68_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_83_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15591_ channels.sample2\[6\] _06397_ _07526_ _03231_ _07527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_139_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13802__A2 _05078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17330_ _00400_ clknet_leaf_86_clk channels.pw1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_14542_ _06460_ _06465_ _06538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11754_ _03813_ _03845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_139_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17261_ _00331_ clknet_leaf_75_clk tt_um_rejunity_sn76489.control_tone_freq\[2\]\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10705_ _02961_ _02777_ _02962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14473_ _06447_ _06469_ _06470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__16752__A1 _03710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15555__A2 _07493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11685_ _03535_ _03771_ _03774_ _03775_ _03776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_16212_ _08083_ _08084_ _08085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13566__A1 _04597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13424_ _05289_ _05377_ _05430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_17192_ _00262_ clknet_leaf_89_clk filters.cutoff_lut\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10636_ _02846_ _02864_ _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_52_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16143_ _07792_ _07881_ _07886_ _08019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_153_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13355_ _05244_ _05361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_134_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10567_ _02816_ _02826_ _02827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_140_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08993__A1 _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12306_ _04311_ _04312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16074_ _07923_ _07952_ _00653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13286_ _05271_ _05291_ _05292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10498_ _02756_ _02757_ _02759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_5_14__f_clk clknet_3_3_0_clk clknet_5_14__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_122_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15025_ _04693_ _05036_ _05042_ _06995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__12215__I _04220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12237_ _04242_ _04243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_114_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12168_ _04173_ _04174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_5_11__f_clk_I clknet_3_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10552__A1 _02535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11119_ filters.sample_filtered\[6\] _03337_ _03338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_36_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16976_ _00055_ clknet_leaf_187_clk channels.accum\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12099_ _01219_ _03551_ _01931_ _04131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_127_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 addr[5] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15927_ _07808_ _07809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_127_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16035__A3 _07914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15858_ _07717_ _07741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12057__A1 _01319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14809_ _06701_ _06794_ _06795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_176_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15261__I _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15789_ _07663_ _07690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_177_3662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_177_3673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17528_ _00598_ clknet_5_6__leaf_clk filters.sample_buff\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16743__A1 _08456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17459_ _00529_ clknet_leaf_4_clk filters.band\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_138_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13557__A1 _05560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14809__A1 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_87_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09715_ _02089_ _02090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_93_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09646_ channels.freq1\[5\] _02011_ _02012_ channels.pw3\[5\] _02032_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__14037__A2 _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_182_Right_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_139_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12795__I _04800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09577_ channels.sus_rel3\[3\] _01963_ _01964_ channels.sus_rel1\[3\] _01965_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_167_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13796__A1 _05794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12599__A2 _04541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08528_ _01027_ _01031_ _01052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_107_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11470_ channels.accum\[1\]\[19\] _03590_ _03619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10421_ _02656_ _02658_ _02654_ _02682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_180_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15120__B _07086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13140_ _04320_ _05145_ _05146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12771__A2 _04776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10352_ _02591_ _02613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08513__I _01008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_1164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13071_ filters.high\[16\] filters.band\[16\] _03185_ _05077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10283_ channels.env_vol\[0\]\[4\] channels.env_vol\[1\]\[4\] channels.ch3_env\[4\]
+ channels.env_vol\[3\]\[4\] _01143_ _01687_ _02544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XTAP_TAPCELL_ROW_76_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12022_ channels.env_counter\[1\]\[4\] _04085_ _04086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11731__C2 channels.atk_dec1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16830_ _03492_ _00925_ _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14276__A2 _06192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11095__B _03314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16761_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[8\] _00873_ _00871_ _00876_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13973_ _04161_ _05973_ _05974_ _00530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_12924_ _04295_ _04929_ _04930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15712_ _05534_ _07633_ _07356_ _07634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16692_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[8\] _08400_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[8\]
+ _08433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__10837__A2 _02890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14028__A2 _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12855_ _04860_ _04861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15643_ channels.sample3\[10\] _07549_ _07575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15776__A2 _07640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11806_ _03890_ _03838_ _03897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13787__A1 _04966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15574_ filters.sample_buff\[5\] _07484_ _07511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12786_ _04311_ _04321_ _04444_ _04791_ _04792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_56_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09455__A2 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14525_ _06520_ _06254_ _06483_ _06521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17313_ _00383_ clknet_leaf_161_clk channels.accum\[1\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11737_ _03801_ _03814_ _03828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_154_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16725__A1 _01800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15528__A2 _07468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_155_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_155_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_127_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17244_ _00314_ clknet_leaf_90_clk filters.sample_filtered\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14456_ _06337_ _06451_ _06452_ _06453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_71_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_172_3570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11668_ channels.sus_rel3\[5\] _01081_ _01281_ channels.sus_rel2\[5\] _03758_ _03759_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_25_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_172_3581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13407_ _05412_ _05411_ _05413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_114_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17175_ _00245_ clknet_leaf_141_clk channels.atk_dec3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_116_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10619_ _02842_ _02877_ _02878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_153_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14387_ _06382_ _06384_ _06385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_11599_ _03689_ _03705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_107_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16126_ _07977_ _07981_ _08002_ _08003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_109_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13338_ _04257_ _04739_ _05344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16057_ _07932_ _07934_ _07935_ _07936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_13269_ _04629_ _05268_ _05275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15008_ _06978_ _06979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10525__A1 _02359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12278__A1 _04252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16959_ _00038_ clknet_leaf_232_clk channels.env_vol\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_154_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_179_3702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09500_ _01890_ _01891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12817__A3 _04784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_179_3713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10828__A2 _03080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_133_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12293__A4 _04296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09431_ _01821_ _01822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_78_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13504__I _04850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09362_ _01762_ _01749_ _01763_ _01764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_23_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16815__I _00914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16716__A1 _08449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09293_ _01717_ _01718_ _01711_ _01719_ _01604_ _01606_ _01720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_145_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09857__C _02103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13950__A1 _04254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11694__I _03784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09164__I _01590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12269__A1 _04274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08568__S0 _00009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10103__I _02365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10970_ filters.filter_step\[0\] _03195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09629_ _02008_ _02010_ _02013_ _02015_ _02016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_74_1265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12640_ _04628_ _04645_ _04635_ _04646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_38_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14430__A2 _05187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12571_ _04354_ _04576_ _04577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_50_clk clknet_5_10__leaf_clk clknet_leaf_50_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_136_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14310_ _06306_ _06307_ _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11522_ _03651_ _03652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15290_ _07246_ _07249_ _07250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_109_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14194__A1 _06105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14241_ _06237_ _06238_ _06239_ _06240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_108_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11453_ channels.accum\[1\]\[12\] _03609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10773__I _02602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09339__I _01741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08948__A1 channels.freq2\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_150_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10404_ _02661_ _02663_ _02665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_150_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08948__B2 channels.freq1\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14172_ _06059_ _06061_ _06172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11384_ channels.accum\[2\]\[8\] _03568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_12_Left_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13123_ _05101_ _05128_ _05129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_103_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10335_ _02591_ _02593_ _02595_ _02596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_108_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13054_ _04922_ _04931_ _05059_ _05060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10266_ _02372_ _02525_ _02526_ _02527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_12005_ _04007_ _04072_ _04073_ _00463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09373__A1 _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10197_ _02454_ _01099_ _02456_ _02457_ _02458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_108_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16813_ _00879_ _00913_ _00914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_75_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16744_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[8\] _00861_ _00863_ _00865_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13956_ _05937_ _05957_ _05958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_88_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12907_ _04833_ _04837_ _04913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_88_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16675_ _06978_ _08419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13887_ _05887_ _05888_ _05889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_157_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15626_ filters.sample_buff\[8\] _07447_ _07523_ _07559_ _07560_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_12838_ _04841_ _04842_ _04843_ _04844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_174_3610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_174_3621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15557_ _07487_ _07480_ _07494_ _07496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_12769_ _04762_ _04774_ _04775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_41_clk clknet_5_3__leaf_clk clknet_leaf_41_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_126_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14508_ _06503_ _06504_ _06505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15488_ _07431_ _07432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_142_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_154_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17227_ _00297_ clknet_leaf_176_clk channels.sample1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_141_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14439_ _06326_ _06327_ _06436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_114_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09287__S1 _01328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09249__I _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12735__A2 _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17158_ _00228_ clknet_leaf_142_clk channels.freq3\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10746__A1 _02676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16109_ _07940_ _07907_ _07986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17089_ _00159_ clknet_leaf_107_clk channels.pw1\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09693__B _02036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09980_ _02245_ _02275_ _02278_ _00233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_122_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10210__A3 channels.pw3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14488__A2 _05560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08931_ _01076_ _01397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_36_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_122_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08862_ _01256_ _01334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08793_ _01265_ _01266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_58_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09414_ _01751_ _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09345_ _01747_ _01748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_48_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_32_clk clknet_5_2__leaf_clk clknet_leaf_32_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_47_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08722__S0 _01152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09276_ _01701_ _01683_ _01705_ _01699_ _00098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_168_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14176__A1 _06168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_95_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09159__I _01304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10737__A1 _02602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_56_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_113_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_179_1300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10120_ channels.ctrl_reg3\[5\] _01074_ _01274_ channels.ctrl_reg2\[5\] _02380_ _02381_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_73_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_99_clk clknet_5_13__leaf_clk clknet_leaf_99_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10051_ _02326_ _02320_ _02327_ _00255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13151__A2 _04896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_175_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09107__A1 _01323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13810_ _05717_ _05738_ _05812_ _05813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_14790_ filters.low\[18\] filters.band\[18\] _06073_ _06778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13741_ _05559_ _05641_ _05745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12662__A1 _04667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10953_ _03174_ _03141_ _03178_ _00306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16460_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[6\] _08255_ _08256_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13672_ _05670_ _05675_ _05676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_167_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10884_ _03126_ _03134_ _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_85_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12623_ _04420_ _04629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15411_ _06822_ _07348_ _07344_ _07352_ _07360_ _07361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_16391_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[4\] _08198_ _08205_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_14_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_23_clk clknet_5_1__leaf_clk clknet_leaf_23_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_14_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_152_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15342_ _07283_ _07296_ _07285_ _07298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_171_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_152_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12965__A2 _04966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12554_ _04528_ _04532_ _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_65_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_81_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11505_ _01740_ _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15273_ _05849_ _05851_ _07233_ _07234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_149_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12485_ _04490_ _04491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_20_Left_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_53_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17012_ _00091_ clknet_leaf_227_clk channels.lfsr\[2\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14224_ _04452_ _05947_ _06223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11436_ _03160_ _01381_ _03598_ _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_130_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09594__A1 channels.atk_dec3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09594__B2 channels.pw3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14155_ _06153_ _06154_ _06155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_21_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11367_ _01311_ _03557_ _01316_ _03558_ _00340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_104_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13106_ _03301_ _04332_ _04783_ _05112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_21_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10318_ _01143_ _02578_ _02579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14086_ _05990_ _06086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11298_ _02314_ _03498_ _03502_ _00327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_167_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13142__A2 _04800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13037_ _04992_ _05016_ _05042_ _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_167_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10249_ _01497_ _02378_ _02510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_28_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_128_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10900__A1 _02366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17776_ _00846_ clknet_leaf_206_clk channels.exp_periods\[1\]\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14988_ _06944_ _06946_ _06959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16727_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[9\] _08454_ _08459_ _08460_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13939_ _04176_ _05796_ _05941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16658_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[1\] _08398_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[1\]
+ _08405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_141_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15609_ filters.sample_buff\[7\] _07543_ _07544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09688__B _02036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16589_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[7\] _08345_ _08339_ _08365_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_146_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_14_clk clknet_5_6__leaf_clk clknet_leaf_14_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_17_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09130_ _01577_ _01578_ _01579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_45_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12956__A2 _04766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09282__B1 _01710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14158__A1 _06142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09061_ _01257_ _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12708__A2 _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10719__A1 channels.sample3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15709__I _07630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09585__A1 channels.atk_dec2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12184__A3 _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10195__A2 _02455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09963_ _02264_ _02266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_60_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_90_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14330__A1 _04446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13133__A2 _04818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08914_ channels.accum\[0\]\[5\] _01360_ _01382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09894_ channels.atk_dec2\[3\] _02211_ _02217_ _02218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_176_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_51_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08845_ _01317_ _01318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08776_ _01072_ _01250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input12_I bus_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09196__S0 _01605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11447__A2 _03605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09328_ _01694_ _01736_ _01737_ _01696_ _00118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_35_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12947__A2 _04482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14149__A1 _06015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09259_ channels.lfsr\[1\]\[15\] _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_105_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12270_ _03180_ _03181_ _03183_ _03298_ _04276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_107_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11221_ filters.sample_filtered\[11\] _03415_ _03433_ _03434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_181_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13372__A2 _05377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11383__A1 _03566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09617__I _01941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11152_ _03368_ _03356_ _03369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10103_ _02365_ _02366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_179_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15960_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[1\] _07841_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_11083_ _03298_ _03207_ _03303_ _03304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10034_ _02314_ _02310_ _02315_ _00250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14911_ _06885_ _06887_ _06888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_249_clk_I clknet_5_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15891_ _07772_ _07773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_145_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16074__A1 _07923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17630_ _00700_ clknet_leaf_213_clk channels.env_vol\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14842_ _06777_ _06824_ _06825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_76_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14624__A2 _04601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_106_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17561_ _00631_ clknet_leaf_30_clk filters.low\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11985_ _04043_ _04056_ _04057_ _00459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14773_ _06762_ _06763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16512_ _08296_ _08299_ _08300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_123_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13724_ _05630_ _05726_ _05727_ _05728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_86_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10936_ channels.sample1\[4\] _03164_ _03169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17492_ _00562_ clknet_leaf_8_clk filters.high\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__16377__A2 _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16443_ _08243_ _08244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13655_ _05568_ _05575_ _05659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_10867_ _03117_ _03118_ _03119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_112_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12606_ _04611_ _04612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_16374_ _08190_ _08191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13586_ _05586_ _05590_ _05591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_38_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10798_ channels.sample3\[6\] _02975_ _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_170_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12537_ _04540_ _04542_ _04543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_15325_ _07035_ _07281_ _07282_ _00574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15888__A1 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[0\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12468_ _04467_ _04471_ _04390_ _04473_ _04474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_83_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15256_ _03422_ _07216_ _07218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14207_ _04737_ _05731_ _06206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11419_ channels.accum\[2\]\[23\] _03556_ _03588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10961__I _03185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15187_ _07128_ _07132_ _07151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_105_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12399_ _04404_ _04405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11374__A1 _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14138_ _06011_ _06019_ _06138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_165_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14069_ _06065_ _06069_ _06070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_33_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_182_3753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input4_I addr[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_182_3775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08630_ channels.lfsr\[3\]\[19\] _01126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08561_ _01077_ _01078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_17759_ _00829_ clknet_leaf_70_clk tt_um_rejunity_sn76489.latch_control_reg\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_178_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08492_ _01016_ _00129_ _01021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10101__A2 _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09113_ channels.accum\[2\]\[22\] _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_165_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09044_ _01436_ _01501_ _01502_ _01503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_60_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_92_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13106__A2 _04332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14303__A1 _06275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09946_ _02174_ _02254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11117__A1 filters.high\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12798__I _04803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09877_ _02157_ _02201_ _02205_ _00203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_5_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08828_ channels.freq3\[0\] _01074_ _01301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10312__S _01142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14606__A2 _06601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_79_Right_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09169__S0 _01141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08759_ channels.exp_counter\[1\]\[4\] _01230_ _01238_ _01101_ _01239_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_68_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10111__I _02371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11770_ channels.env_counter\[0\]\[5\] channels.env_counter\[1\]\[5\] channels.env_counter\[2\]\[5\]
+ channels.env_counter\[3\]\[5\] _01152_ _01171_ _03861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_36_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10721_ _02972_ _02977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_55_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13440_ _04596_ _05446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10652_ _02644_ _02775_ _02910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08516__I _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09797__A1 _02131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13593__A2 _05596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13371_ _05376_ _05293_ _05377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_64_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16733__I _08463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10583_ _02838_ _02841_ _02842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_91_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12322_ _04319_ _04327_ _04328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_88_Right_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15110_ _07069_ _07072_ _07076_ _07077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_16090_ _07963_ _07967_ _07968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_106_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16531__A2 _08315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_173_clk_I clknet_5_24__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09549__A1 channels.sus_rel2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15041_ _07008_ _06996_ _07009_ _07010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_160_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09549__B2 channels.freq3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12253_ _04258_ _04259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__11356__A1 _03529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09347__I _01062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_53_clk_I clknet_5_10__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11204_ _03417_ _03407_ _03418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_31_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11098__B _03317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12184_ _03239_ _03203_ _04189_ _03343_ _04190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_147_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15098__A2 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08772__A2 _01245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11135_ filters.sample_filtered\[7\] _03352_ _03353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_43_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_188_clk_I clknet_5_19__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16992_ _00071_ clknet_leaf_155_clk channels.accum\[0\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15943_ _07813_ _07825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_11066_ _03287_ _03288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_leaf_68_clk_I clknet_5_11__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09721__A1 channels.pw1\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10017_ channels.atk_dec3\[4\] _02302_ _02303_ _02304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_125_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_97_Right_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_160_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_160_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15874_ _07755_ tt_um_rejunity_sn76489.chan\[2\].attenuation.in _07756_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_111_clk_I clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17613_ _00683_ clknet_leaf_135_clk channels.env_counter\[3\]\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14825_ _06804_ _06809_ _06810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_116_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15270__A2 _07230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17544_ _00614_ clknet_leaf_0_clk filters.low\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_175_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14756_ _05544_ _06746_ _06747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11968_ _04006_ _04043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13707_ _05619_ _05709_ _05710_ _05711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17475_ _00545_ clknet_leaf_244_clk filters.band\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10919_ _03154_ _03122_ _03158_ _00292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14687_ _06664_ _06667_ _06681_ _06682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_11899_ _03960_ _03981_ _03982_ _00448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_156_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16426_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[13\] _08223_ _08230_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13638_ _05553_ _05642_ _05643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_6_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_172_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13584__A2 _05588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16357_ channels.ch3_env\[1\] _08179_ _08181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14781__A1 _06769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13569_ _05572_ _05573_ _05574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_4_Left_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11595__A1 channels.pw3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15308_ _07265_ _07266_ _07086_ _07267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16288_ _02354_ _03741_ _00678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_164_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13336__A2 _04860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15239_ _07198_ _07199_ _07200_ _07201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_140_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16286__A1 _02103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09800_ _02141_ _02151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09960__A1 _02242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08763__A2 _01090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13639__A3 _05643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09731_ _02102_ _02103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_163_Right_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12847__A1 _04476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09712__A1 _01819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09662_ _02043_ _02044_ _02045_ _02046_ _02047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_94_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08613_ _01117_ _00023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09593_ channels.pw2\[3\] _01847_ _01900_ channels.atk_dec1\[3\] _01981_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_55_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08544_ _00132_ _01061_ _01044_ _00008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10086__A1 net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08475_ _01004_ _01005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_49_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09779__A1 _01807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09027_ _01449_ _01486_ _01487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09929_ _02240_ _02235_ _02241_ _00219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_130_Right_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_142_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12940_ _04945_ _04946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_12871_ _04828_ _04838_ _04877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_87_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14610_ _06503_ _06604_ _06605_ _06606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11822_ _03904_ _03908_ _03910_ _03912_ _03913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_96_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_83_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15590_ _03342_ _07513_ _07525_ _06177_ _07526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_83_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10077__A1 _02326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11753_ _03841_ _03843_ _03844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_28_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14541_ _06535_ _06536_ _06537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11813__A2 _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13152__I _04366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09482__A3 _01865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10704_ _02657_ _02961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17260_ _00330_ clknet_leaf_74_clk tt_um_rejunity_sn76489.control_tone_freq\[2\]\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09219__B1 _01657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14472_ _06450_ _06468_ _06469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11684_ _03536_ _03535_ _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_154_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16211_ _07960_ _08014_ _07988_ _07786_ _08084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_52_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13566__A2 _05570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10635_ _02846_ _02864_ _02893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13423_ _05427_ _05428_ _05429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_125_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17191_ _00261_ clknet_leaf_89_clk filters.cutoff_lut\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_36_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11577__A1 channels.freq3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16142_ _07801_ _07786_ _07800_ _07794_ _08018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_23_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13354_ _05278_ _05282_ _05359_ _05360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_3_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10566_ _02819_ _02825_ _02826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__16504__A2 _08289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12305_ _03199_ _04216_ _04311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_87_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16073_ spi_dac_i.spi_dat_buff_1\[3\] _07924_ _07951_ _07952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13285_ _05274_ _05290_ _05291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10497_ _02756_ _02757_ _02758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_122_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13869__A3 _05849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12236_ _04241_ _04242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15024_ _05016_ _06994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_122_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16268__A1 filters.sample_buff\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09942__A1 _02250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10016__I _02293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12167_ filters.res_lut\[1\] _04167_ _04173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09805__I _02154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10552__A2 _02500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11118_ _03334_ _03336_ _03337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_12098_ _04130_ _00499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12829__A1 _04316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16975_ _00054_ clknet_leaf_193_clk channels.ring_outs\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15926_ tt_um_rejunity_sn76489.chan\[3\].attenuation.in _07808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_11049_ _03271_ _03272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput7 bus_cyc net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11501__A1 channels.freq1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15857_ _07730_ _07739_ _07740_ _00648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_59_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14046__A3 _05721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14808_ filters.low\[20\] filters.band\[20\] _03472_ _06794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_87_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15788_ _07688_ _07689_ _00630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_146_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10068__A1 _02299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_177_3663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17527_ _00597_ clknet_leaf_19_clk filters.sample_buff\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14739_ _03456_ _03222_ _06730_ _06731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_177_3674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_172_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_145_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17458_ _00528_ clknet_leaf_1_clk filters.band\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_138_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16409_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[9\] _08209_ _08218_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17389_ _00459_ clknet_leaf_148_clk channels.env_counter\[2\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11568__A1 _03662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14822__S _06073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11310__I _02184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12368__I0 filters.cutoff_lut\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09933__A1 _02242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09714_ _02088_ _01891_ _02089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_179_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09645_ channels.ch3_env\[5\] _02009_ _01948_ channels.atk_dec1\[5\] _02031_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09576_ _01898_ _01964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_132_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08527_ _01051_ _00130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_171_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_20__f_clk clknet_3_5_0_clk clknet_5_20__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_61_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10420_ _02675_ _02679_ _02680_ _02681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_0_45_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09621__B1 _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10351_ _02585_ _02596_ _02612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_182_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13070_ _04175_ _05075_ _05076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10282_ _02538_ _02540_ _02542_ _02543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_13_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_76_Left_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12021_ _04077_ _04085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_76_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13720__A2 _05723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11731__B2 channels.atk_dec2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_5_3__f_clk_I clknet_3_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16760_ _08456_ _00868_ _00875_ _00809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13484__A1 _05484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13972_ filters.band\[4\] _05540_ _05541_ _05974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09152__A2 _01592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15711_ _07630_ _07633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12923_ _04491_ _04929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_77_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16691_ _08431_ _08432_ _00790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_88_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15225__A2 _07187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15642_ filters.sample_buff\[9\] _07568_ _07574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12854_ filters.high\[14\] filters.band\[14\] _04710_ _04860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_158_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_85_Left_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11805_ _03881_ _03882_ _03883_ _03895_ _03896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_139_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13787__A2 _04447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15573_ _07498_ _07510_ _00594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_115_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12785_ _04783_ _04791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_173_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17312_ _00382_ clknet_leaf_157_clk channels.accum\[1\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14524_ _06484_ _06520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_113_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11736_ _03825_ _03826_ _03827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_127_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17243_ _00313_ clknet_leaf_91_clk filters.sample_filtered\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14736__A1 _06403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14455_ _06334_ _06344_ _06452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14706__I _06688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11667_ channels.sus_rel1\[5\] _01294_ _03758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_126_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_172_3571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_172_3582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13406_ _05394_ _05395_ _05397_ _05412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_52_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17174_ _00244_ clknet_leaf_118_clk channels.atk_dec3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10618_ _02844_ _02876_ _02877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_148_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11598_ _03695_ _03704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14386_ _05563_ _06383_ _06384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16125_ _07985_ _08001_ _08002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_84_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10549_ _02800_ _02808_ _02809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13337_ net57 _04711_ _05343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_94_Left_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16056_ _07774_ _07778_ _07780_ _07935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13268_ _05168_ _05272_ _05273_ _05274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_122_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15007_ _03940_ _06978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12219_ _04224_ _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13199_ _05151_ _05205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10525__A2 _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16661__A1 _08333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15464__A2 _06717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16796__C _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16958_ _00037_ clknet_5_16__leaf_clk channels.env_vol\[3\]\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_179_3703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15909_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[2\] _07790_ _07791_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_179_3714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16889_ _01193_ _00938_ _00972_ _00841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_200_clk clknet_5_23__leaf_clk clknet_leaf_200_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09430_ _01102_ _01821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_78_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09361_ _01752_ _01763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_87_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09292_ channels.lfsr\[3\]\[21\] _01719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_129_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_160_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13950__A2 _05185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09906__A1 _02160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08590__B1 _01105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08568__S1 _00010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15207__A2 _07146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09628_ filters.lp _02014_ _01964_ channels.sus_rel1\[4\] _02015_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_168_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14966__A1 _05647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09559_ _01900_ _01948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_66_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_136_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12570_ _04575_ _04576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11521_ _02333_ _03651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_135_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_81_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11452_ _03600_ _01459_ _03608_ _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14240_ filters.band\[27\] _04599_ _06239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14194__A2 _06135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10403_ _02661_ _02663_ _02664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_78_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14171_ _06059_ _06061_ _06171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_78_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_150_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11383_ _03566_ _01406_ _03567_ _00347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_150_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10334_ _02509_ _02528_ _02594_ _02595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_13122_ _05115_ _05127_ _05128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_103_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13053_ _04917_ _04921_ _05059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__16891__A1 _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10265_ _01497_ _02382_ _02526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_178_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12004_ channels.env_counter\[2\]\[14\] _04012_ _04073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09355__I _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11704__B2 channels.atk_dec2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10196_ channels.pw1\[2\] _02430_ _02457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16812_ _08461_ _08442_ _00880_ _00893_ _01817_ _01811_ _00913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai33_1
XANTENNA__15446__A2 _06934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16743_ _08456_ _08464_ _00864_ _00803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13955_ _05940_ _05956_ _05957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_159_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12906_ _04833_ _04837_ _04912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16674_ _08356_ _08418_ _00787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13886_ _05789_ _05810_ _05888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_76_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15625_ _07557_ _07558_ _07559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10691__A1 _02686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14957__A1 _06921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12837_ _04732_ _04736_ _04843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_174_3611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_174_3622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15556_ _07487_ _07480_ _07494_ _07495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_16_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12768_ _04772_ _04773_ _04774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14507_ _06298_ _06400_ _06504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11719_ _03788_ _03809_ _03810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_16_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15487_ _07416_ _07428_ _07430_ _07431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_12699_ _04476_ _04705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_182_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17226_ _00296_ clknet_leaf_176_clk channels.sample1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput10 bus_in[2] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_14438_ _06433_ _06434_ _06435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_71_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12196__A1 _03288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_249_clk clknet_5_1__leaf_clk clknet_leaf_249_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_109_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17157_ _00227_ clknet_leaf_142_clk channels.freq3\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14369_ _06361_ _06366_ _06367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__15695__C _07269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10746__A2 _02872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16108_ _07982_ _07984_ _07985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_17088_ _00158_ clknet_leaf_112_clk channels.pw1\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_110_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11795__I _01149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16039_ _07916_ _07918_ _07919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08930_ _01389_ _01390_ _01396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_23_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_36_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08861_ _01323_ _01331_ _01332_ _01333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_97_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16600__B _08318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15437__A2 _06765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08792_ _01096_ _01265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09116__A2 _01566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09413_ _01806_ _01807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_149_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15730__I _07355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09344_ _01746_ _01747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09275_ _01702_ _01703_ _01700_ _01704_ _01144_ _01158_ _01705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__08722__S1 _01168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12187__A1 _03350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13923__A2 _04818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_56_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13687__A1 _04400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10050_ channels.sus_rel3\[6\] _02321_ _02322_ _02327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13439__A1 _04561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13740_ _05559_ _05641_ _05744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_138_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10952_ channels.sample1\[11\] _01261_ _03178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16928__A2 _00993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13671_ _05673_ _05674_ _05675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_35_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10883_ _03127_ _03133_ _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__15640__I _06978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15410_ _07351_ _07360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_12622_ _04354_ _04628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_94_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16390_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[3\] _08201_ _08204_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_159_Left_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_152_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10784__I _02676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15341_ _07283_ _07296_ _07297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12553_ _04549_ _04545_ _04546_ _04559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_108_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11504_ _02328_ _03632_ _03638_ _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_15272_ _07232_ _07233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_12484_ _04489_ _04490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12178__A1 filters.res_lut\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17011_ _00090_ clknet_leaf_227_clk channels.lfsr\[2\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14223_ _04326_ _05501_ _06222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11435_ channels.accum\[1\]\[5\] _03593_ _03598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12705__S _04710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_130_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14154_ _04230_ _05588_ _06154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11366_ _01084_ _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_132_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10317_ channels.ch3_env\[5\] _02578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13105_ net64 _04196_ _04779_ _05111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11297_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[1\] _03500_ _03485_ _03502_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14085_ _05997_ _06083_ _06084_ _06085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13678__A1 _05594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_168_Left_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_167_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10248_ _02508_ _02509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13036_ _05039_ _05040_ _05041_ _05042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_167_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11153__A2 _03352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10179_ _02426_ _02428_ channels.pw3\[4\] _02440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_128_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10900__A2 _02880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16092__A2 _07942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17775_ _00845_ clknet_leaf_204_clk channels.exp_periods\[1\]\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15036__B _06979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14987_ _06935_ _06950_ _06957_ _06958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_178_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16726_ _08450_ _08459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_152_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13938_ _05816_ _05824_ _05939_ _05940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_77_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10664__A1 _01085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16657_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[2\] _08398_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[2\]
+ _08404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13869_ _05747_ _05870_ _05849_ _05871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XPHY_EDGE_ROW_177_Left_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_141_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15608_ _07541_ _07542_ _07543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_16588_ _08333_ _08362_ _08363_ _08364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_173_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15539_ filters.sample_buff\[2\] _07478_ _07479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_45_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09282__B2 _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09060_ channels.accum\[0\]\[16\] _01517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17209_ _00279_ clknet_leaf_94_clk channels.sample3\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09034__A1 channels.freq2\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09034__B2 channels.freq1\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_38_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10195__A3 channels.pw3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09962_ _02264_ _02265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08913_ _01349_ _01380_ _01381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09893_ _02216_ _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_51_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08844_ _01253_ _01317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_58_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_100_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08775_ _01248_ _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14094__A1 _05446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09196__S1 _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08848__A1 _01070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14397__A2 _06394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09327_ _01730_ _01737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14149__A2 _06016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15346__A1 _06983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09258_ channels.lfsr\[0\]\[15\] _01691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_32_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09189_ _01629_ _01630_ _01621_ _01631_ _01141_ _01155_ _01632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_160_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_177_Right_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11220_ _03432_ _03419_ _03433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_31_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12580__A1 _04574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11151_ _03353_ _03368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_105_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10102_ _02364_ _02365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11082_ filters.low\[4\] _03217_ _03302_ _03207_ _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_101_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11135__A2 _03352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10033_ channels.sus_rel3\[1\] _02311_ _02312_ _02315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14910_ _06874_ _06878_ _06886_ _06887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15890_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[2\] _07765_ _07772_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_145_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14841_ _06822_ _03473_ _06823_ _06824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15821__A2 _07631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17560_ _00630_ clknet_leaf_29_clk filters.low\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_106_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08839__A1 _01308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14772_ _03733_ _06762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_106_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11984_ channels.env_counter\[2\]\[10\] _04048_ _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13832__A1 _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16511_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[6\] _08269_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[6\]
+ _08299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_123_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13723_ _05631_ _05632_ _05727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_86_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17491_ _00561_ clknet_leaf_243_clk filters.high\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10935_ _01320_ _03168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_168_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16442_ _08242_ _08243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13654_ net35 net40 _05531_ _05643_ _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_10866_ _03094_ _03098_ _03118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_38_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12605_ _04577_ _04580_ _04611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_16373_ tt_um_rejunity_sn76489.noise\[0\].gen.signal_edge.previous_signal_state_0
+ _02349_ _08190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_27_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13585_ _05587_ _05589_ _05590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_38_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10797_ _03018_ _03051_ _03052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_53_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10949__A2 _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15324_ filters.high\[16\] _07062_ _07223_ _07282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12536_ _04165_ _04541_ _04542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_82_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09016__A1 _01468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15255_ filters.low\[12\] _07216_ _07217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_12467_ _04279_ _04473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13899__A1 _05813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09808__I _01813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_144_Right_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_14206_ _04750_ _05625_ _06205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_169_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11418_ _01564_ _03581_ _01568_ _03582_ _00362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_111_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15186_ _07128_ _07132_ _07150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12398_ _03398_ _04403_ _04404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_10_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14137_ _06014_ _06018_ _06137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11349_ _03535_ _03542_ _03543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_33_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14068_ _03314_ _06067_ _06068_ _06069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_20_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15545__I _07446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13019_ _04462_ _05006_ _05025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_182_3776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_182_3787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__16065__A2 _07914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08560_ _01076_ _01077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17758_ _00828_ clknet_leaf_81_clk tt_um_rejunity_sn76489.noise\[0\].gen.restart_noise
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_16709_ _08445_ _08447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08491_ _01020_ _00129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_175_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17689_ _00759_ clknet_leaf_63_clk tt_um_rejunity_sn76489.chan\[1\].attenuation.in
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_175_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_5_1__f_clk clknet_3_0_0_clk clknet_5_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_58_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_1300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11313__I _02187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09112_ channels.accum\[1\]\[22\] _01563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_165_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09043_ _01491_ _01485_ _01500_ _01502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_44_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14000__A1 _05950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_111_Right_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__16828__A1 _00923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09945_ _02252_ _02247_ _02253_ _00223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13106__A3 _04783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14303__A2 _06277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09876_ channels.ctrl_reg2\[6\] _02202_ _02199_ _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_5_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08827_ _01299_ _01300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14067__A1 _03310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15803__A2 _07631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09169__S1 _01155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08758_ _01217_ _01237_ _01238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_174_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08689_ _01172_ _01173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_138_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10720_ _02882_ _02973_ _02976_ _00275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_165_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15567__A1 filters.sample_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12319__I _04324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10651_ _02657_ _02622_ _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_81_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13370_ _05375_ _05295_ _05376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10582_ _02839_ _02819_ _02840_ _02841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_36_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13593__A3 _05597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12396__A4 filters.high\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16235__B _07741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12321_ _04322_ _04326_ _04327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_133_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15040_ _05969_ _06993_ _07009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_142_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12252_ _04257_ _04258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_146_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11356__A2 _03531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11203_ _03404_ _03417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12183_ _04188_ _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_147_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11134_ _03343_ _03344_ _03351_ _03352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_16991_ _00070_ clknet_5_28__leaf_clk channels.accum\[0\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12305__A1 _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15942_ _07820_ _07823_ _07824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11065_ net63 _03287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10016_ _02293_ _02303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_125_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17495__CLK clknet_5_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15873_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[2\] _07755_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_160_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_160_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17612_ _00682_ clknet_leaf_129_clk channels.env_counter\[3\]\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14824_ _06806_ _06808_ _06809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_157_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13805__A1 _05803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12608__A2 _04171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17543_ _00613_ clknet_leaf_243_clk filters.low\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14755_ _06742_ _06745_ _06746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11967_ _04027_ _04041_ _04042_ _00456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13706_ _05620_ _05621_ _05710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_17474_ _00544_ clknet_leaf_244_clk filters.band\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10918_ channels.sample2\[9\] _03156_ _03158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14686_ _06668_ _06674_ _06680_ _06681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_54_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11898_ channels.env_vol\[0\]\[7\] _03965_ _03982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16425_ _08228_ _08229_ _08222_ _00727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13637_ _05555_ _05559_ _05641_ _05642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_6_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10849_ _03099_ _03101_ _03102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_67_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10177__C _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16356_ _03743_ _08177_ _08180_ _00707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_172_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13568_ _04764_ _05570_ _05573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15307_ _07246_ _07249_ _07256_ _07266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_12519_ _04266_ _04525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_125_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16287_ _03738_ _03740_ _00677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13499_ _05504_ _05505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15238_ _07176_ _07191_ _07200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09096__S0 _01138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15169_ filters.low\[9\] _07133_ _07134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__16286__A2 _07838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09730_ _02101_ _02102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09661_ channels.pw1\[6\] _02003_ _02004_ channels.ctrl_reg1\[6\] _02046_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__14049__A1 _04372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_105_Left_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_173_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08612_ channels.lfsr\[3\]\[10\] _01117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09592_ channels.ctrl_reg2\[3\] _01974_ _01882_ channels.ctrl_reg3\[3\] _01979_ _01980_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_55_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08543_ _00131_ _01033_ _01061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_148_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_233_clk_I clknet_5_17__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10086__A2 _02351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08474_ _01002_ _01003_ _01004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_46_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_148_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_114_Left_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_116_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_248_clk_I clknet_5_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09026_ _01484_ _01485_ _01486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11199__B _03412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09087__S0 _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11338__A2 _03531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12535__A1 filters.res_lut\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09400__A1 _01757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09928_ channels.sus_rel2\[6\] _02236_ _02232_ _02241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09183__I _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09859_ _02193_ _02194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_176_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12870_ _04840_ _04869_ _04875_ _04876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_38_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11821_ _03906_ _03847_ _03911_ _03912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__09467__A1 channels.freq1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13263__A2 _05268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09467__B2 channels.ctrl_reg1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14460__A1 _06456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11274__A1 _02088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14540_ _06447_ _06469_ _06536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11752_ channels.env_counter\[0\]\[9\] channels.env_counter\[1\]\[9\] channels.env_counter\[2\]\[9\]
+ channels.env_counter\[3\]\[9\] _03832_ _03842_ _03843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_56_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10703_ _02710_ _02873_ _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14471_ _06453_ _06467_ _06468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_37_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11683_ _03748_ _02752_ _03766_ _03039_ _03774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_16210_ _07933_ _07777_ _07930_ _07792_ _08083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_138_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_126_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13422_ _05405_ _05415_ _05417_ _05420_ _05428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_17190_ _00260_ clknet_leaf_78_clk filters.cutoff_lut\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10634_ _02889_ _02891_ _02892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_153_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16141_ _07933_ _08015_ _08016_ _07893_ _08017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_36_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13353_ _04500_ _05092_ _05283_ _05359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_106_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10565_ _02607_ _02824_ _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_118_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12304_ _04213_ _04306_ _04310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_16072_ _07948_ _07949_ _07950_ _07869_ _07951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__13318__A3 _05220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15712__A1 _05534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13284_ _05284_ _05290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_51_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10496_ _02536_ _02554_ _02757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09078__S0 _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12526__A1 _04233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15023_ _06984_ _06992_ _06993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12235_ _04240_ _04241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_20_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12166_ _04165_ _04171_ _04172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__14279__A1 _06275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11117_ filters.high\[6\] _03335_ _03336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12097_ _03554_ channels.adsr_state\[2\]\[1\] _04128_ _04130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12829__A2 _04480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16974_ _00053_ clknet_leaf_191_clk channels.exp_counter\[2\]\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15925_ _07806_ _07807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_11048_ _03270_ _03271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput8 bus_in[0] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_127_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10032__I _02184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15856_ _01822_ _07740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_87_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14807_ _06792_ _06793_ _00545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_15787_ filters.low\[20\] _07682_ _07684_ _07689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_176_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12999_ _05004_ _05005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17526_ _00596_ clknet_leaf_19_clk filters.sample_buff\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14738_ _03455_ _06397_ _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_177_3664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_177_3675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_20__f_clk_I clknet_3_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17457_ _00527_ clknet_leaf_4_clk filters.band\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14669_ _06332_ _06086_ _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16408_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[8\] _08212_ _08217_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_138_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17388_ _00458_ clknet_leaf_149_clk channels.env_counter\[2\]\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13557__A3 _05451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16339_ channels.env_vol\[1\]\[7\] _08166_ _08170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14174__I _06173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13309__A3 _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14506__A2 _06399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12517__A1 _03333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_87_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09713_ _01780_ _02088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09697__A1 _01757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09644_ filters.res_filt\[5\] _02007_ _01939_ _02029_ _02030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_97_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_179_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_172_clk_I clknet_5_24__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09575_ _01943_ _01963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_65_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13245__A2 _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14442__A1 _04355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_167_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08526_ _01043_ _01040_ _01051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_52_clk_I clknet_5_10__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_122_Left_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_187_clk_I clknet_5_19__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_67_clk_I clknet_5_11__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09621__B2 channels.sample3\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_110_clk_I clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10350_ _02606_ _02609_ _02610_ _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_182_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09009_ _01469_ _01470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_42_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10281_ _01482_ _02541_ _02542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10117__I _02377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15170__A2 _07122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12020_ _04074_ _04084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_143_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_131_Left_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_178_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_125_clk_I clknet_5_27__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13971_ _05869_ _05972_ _05973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09688__A1 net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13484__A2 _05489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15710_ _07631_ _07632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_12922_ _04487_ _04927_ _04928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16690_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[7\] _08289_ _01753_ _08432_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_154_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15641_ _07561_ _07572_ _07573_ _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_115_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14028__A4 _06027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12853_ _04174_ _04858_ _04859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_150_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11804_ _03860_ _03861_ _03889_ _03894_ _03895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_15572_ filters.sample_buff\[4\] _07461_ _07451_ _07509_ _07510_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_90_1261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_140_Left_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12784_ _04720_ _04788_ _04789_ _04790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_96_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17311_ _00381_ clknet_leaf_192_clk channels.accum\[1\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14523_ _06471_ _06488_ _06518_ _06519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11735_ _03813_ _03823_ _03826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_25_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17242_ _00312_ clknet_leaf_11_clk filters.sample_filtered\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_155_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14454_ _06342_ _06451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_11666_ _03756_ _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_148_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15311__C _07269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_172_3572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13405_ _04935_ _04950_ _05410_ _05411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_172_3583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17173_ _00243_ clknet_leaf_125_clk channels.atk_dec3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_154_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10617_ _02846_ _02864_ _02875_ _02876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_64_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14385_ _06261_ _06383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_141_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11597_ _03695_ _03703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09088__I _01541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16124_ _07987_ _08000_ _08001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13336_ _04227_ _04860_ _05342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10548_ _02803_ _02806_ _02807_ _02808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_133_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16055_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[2\] _07933_ _07891_
+ _07934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_122_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13267_ _05171_ _05190_ _05273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__15161__A2 _01977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10479_ _02612_ _02650_ _02740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15006_ _06958_ _06975_ _06976_ _06977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12218_ _03311_ _03379_ _03313_ filters.high\[1\] _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XANTENNA__13711__A3 _05714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13198_ _05142_ _05147_ _05204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12149_ _04156_ _00524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09679__A1 channels.freq2\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16957_ _00036_ clknet_leaf_233_clk channels.env_vol\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09679__B2 channels.freq1\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12278__A3 _04283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15908_ _07787_ _07790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11486__A1 channels.freq1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_179_3704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16888_ _00939_ _00971_ _00972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_154_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15839_ spi_dac_i.counter\[4\] _07724_ _07725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13073__I _05078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09360_ _01761_ _01762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_176_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12986__A1 _04952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17509_ _00579_ clknet_leaf_246_clk filters.high\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09291_ channels.lfsr\[1\]\[21\] _01718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_170_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10461__A2 _02721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_83_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_172_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09603__A1 channels.sus_rel3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09603__B2 channels.freq1\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_162_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10213__A2 _02473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09726__I net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13163__A1 _05121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12910__A1 _04855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12152__I _01093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08590__A1 _01086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08590__B2 channels.ring_outs\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15207__A3 _07149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09627_ _01791_ _02014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_69_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09558_ _01935_ _01938_ _01946_ _01947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__16508__B _08292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08509_ _01016_ _01036_ _01037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09489_ _01879_ _01880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11520_ _03641_ _03650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14718__A2 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12729__A1 _04258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11451_ channels.accum\[1\]\[11\] _03605_ _03608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10402_ _02662_ _02645_ _02663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_150_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10204__A2 channels.pw1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14170_ _06169_ _06170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_78_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_150_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11382_ channels.accum\[2\]\[7\] _03559_ _03567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_150_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13121_ _05117_ _05121_ _05126_ _05127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_10333_ _02544_ _02594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13154__A1 _03348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13052_ _05053_ _05057_ _05058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_111_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10264_ _01482_ _02378_ _02525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__16891__A2 _00973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12003_ _03925_ _04070_ _04071_ _04072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10195_ _01582_ _02455_ channels.pw3\[2\] _02456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_100_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16811_ _08456_ _00906_ _00912_ _00910_ _00823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_108_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16742_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[7\] _00861_ _00863_ _00864_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13954_ _05946_ _05955_ _05956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_117_1308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12905_ _04908_ _04909_ _04910_ _04911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16673_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[4\] _08347_ _08416_ _08417_
+ _08418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_13885_ _05792_ _05809_ _05887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_53_1307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_194_clk clknet_5_23__leaf_clk clknet_leaf_194_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_159_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11406__I _01240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15624_ _07548_ _07546_ _07556_ _07558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_124_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12836_ _04744_ _04842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10691__A2 _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_174_3612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15555_ filters.sample_buff\[3\] _07493_ _07494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_5_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11850__B _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12767_ _04748_ _04761_ _04773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_33_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14506_ _06396_ _06399_ _06503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11718_ channels.atk_dec1\[2\] channels.sus_rel1\[2\] _03784_ _03809_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_12_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15486_ _07416_ _06768_ _07429_ _07428_ _07430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_56_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12698_ _04703_ _04180_ _04704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14437_ _06332_ _05671_ _06341_ _06434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_17225_ _00295_ clknet_leaf_170_clk channels.sample1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xinput11 bus_in[3] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_11649_ _01583_ _03739_ _03741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_154_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09597__B1 _01862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17156_ _00226_ clknet_leaf_141_clk channels.freq3\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14368_ _06362_ _06365_ _06366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09974__C _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16107_ _07983_ _07875_ _07955_ _07984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_123_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13319_ _05218_ _05221_ _05324_ _05325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_17087_ _00157_ clknet_leaf_107_clk channels.pw1\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_161_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14299_ _06180_ _06286_ _06297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16038_ _07845_ _07864_ _07917_ _07918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_110_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13068__I _04926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08860_ _01324_ _01330_ _01332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_36_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08791_ _01263_ _01264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_35_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14645__A1 _06472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_185_clk clknet_5_22__leaf_clk clknet_leaf_185_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_176_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09412_ _01805_ _01806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_149_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12959__A1 _04512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09343_ _01745_ _01746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_164_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09824__A1 _02112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_158_Right_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_117_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09274_ channels.lfsr\[3\]\[18\] _01704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_62_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_95_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11934__A2 _03874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_73_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13687__A2 _05690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08989_ channels.freq3\[11\] _01079_ _01451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12610__I _04578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10951_ _03174_ _03136_ _03177_ _00305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10122__A1 channels.ctrl_reg3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_176_clk clknet_5_18__leaf_clk clknet_leaf_176_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13670_ _04211_ _05671_ _05674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10882_ _03130_ _03129_ _03132_ _03133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_156_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16238__B _08098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12621_ _04612_ _04625_ _04626_ _04627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_149_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13441__I _05260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_125_Right_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15340_ _07295_ _06294_ _07296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_54_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12552_ _04556_ _04557_ _04558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_152_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14981__B _06952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11503_ channels.freq1\[7\] _03633_ _03634_ _03638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15271_ filters.low\[13\] _07231_ _07232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_149_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12483_ _03413_ _04488_ _04489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_136_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17010_ _00089_ clknet_leaf_227_clk channels.lfsr\[2\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14222_ _06118_ _06119_ _06220_ _06221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_22_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11434_ _03597_ _03591_ _01372_ _03592_ _00368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10189__A1 _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_145_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14153_ _06151_ _06152_ _06153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_100_clk clknet_5_13__leaf_clk clknet_leaf_100_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_21_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11365_ _03556_ _03557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09366__I _01766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13104_ _03315_ _04163_ _04443_ _05110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_10316_ _02524_ _02569_ _02576_ _02577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_104_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14084_ _06000_ _06057_ _06084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11296_ _03489_ _03498_ _03501_ _02273_ _00326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_46_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16701__B _08318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13035_ _05017_ _05029_ _05038_ _05041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10247_ _02507_ _02508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_167_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12886__B1 _04378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12350__A2 _04355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10178_ channels.pw1\[4\] _02439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_128_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17774_ _00844_ clknet_leaf_202_clk channels.exp_periods\[1\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14986_ _06938_ _06949_ _06957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16725_ _01800_ _08447_ _08458_ _00798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10113__A1 channels.ctrl_reg3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13937_ _05818_ _05938_ _05823_ _05939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_57_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10040__I _02149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16656_ _08356_ _08403_ _00784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13868_ _05531_ _05643_ _05870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_159_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_141_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12676__B _04681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12819_ _04824_ _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_69_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10975__I _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15607_ channels.sample1\[7\] _03427_ _07542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16587_ _08358_ _08361_ _08363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09806__A1 channels.sus_rel1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13799_ _04694_ _05800_ _05091_ _05079_ _05802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_8_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11613__A1 channels.pw2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10416__A2 _02676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15538_ _07476_ _07477_ _07478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_121_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15469_ _07312_ _07413_ _07414_ _00586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_142_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17208_ _00278_ clknet_5_24__leaf_clk channels.sample3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17139_ _00209_ clknet_leaf_127_clk channels.atk_dec2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__15107__A2 channels.sample2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09961_ _01781_ _01842_ _02264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__16855__A2 _03128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08912_ _01374_ _01379_ _01380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_110_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09892_ _02174_ _02216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_176_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11775__S1 _01167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08843_ _01300_ _01315_ _01316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08774_ channels.clk_div\[2\] _01248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_158_clk clknet_5_28__leaf_clk clknet_leaf_158_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08848__A2 _01319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13841__A2 _05813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15741__I _07639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15594__A2 _07529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09326_ _01728_ _01736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11604__A1 channels.pw3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12801__B1 _04806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09257_ channels.lfsr\[2\]\[16\] _01690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_35_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_32_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09188_ channels.lfsr\[3\]\[5\] _01631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_90_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11150_ filters.sample_filtered\[8\] _03366_ _03367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__16521__B _08252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10101_ _01070_ _02363_ _02364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10125__I _02385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11081_ _03301_ _03302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_101_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10032_ _02184_ _02314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_179_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17055__D _00125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14840_ filters.band\[23\] _06755_ _06823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_162_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14771_ _06760_ _06761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_106_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11983_ _04044_ _04055_ _04056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_149_clk clknet_5_31__leaf_clk clknet_leaf_149_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_106_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13832__A2 _04818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16510_ _08265_ _08298_ _00743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13722_ _05631_ _05632_ _05726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_123_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10934_ _03162_ _02932_ _03167_ _00298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_123_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17490_ _00560_ clknet_leaf_13_clk filters.high\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_86_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_169_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16441_ _08241_ _08242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13653_ _05654_ _05655_ _05656_ _05657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_39_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10865_ _03091_ _03093_ _03117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13596__A1 _05584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12604_ _04592_ _04608_ _04609_ _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_156_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16372_ _03981_ _08184_ _08189_ _00714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_155_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13584_ _04400_ _05588_ _05589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10796_ _03049_ _03050_ _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_82_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15323_ _07277_ _07280_ _07281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_12535_ filters.res_lut\[2\] _04169_ _04541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_109_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15254_ _07206_ _07210_ _07215_ _07216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_151_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12466_ _04467_ _04468_ _04469_ _04471_ _04472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__09016__A2 _01470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13899__A2 _05843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14205_ _06202_ _06203_ _06204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_124_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11417_ _03578_ _01559_ _03587_ _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_169_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15185_ _07147_ _07148_ _07149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_12397_ _04402_ _04403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_50_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14136_ _06105_ _06135_ _06136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__12571__A2 _04576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11348_ _03538_ _03541_ _03542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__10582__A1 _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10035__I _02187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14067_ _03310_ _03377_ _06068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11279_ filters.cutoff_lut\[7\] _03483_ _03485_ _03487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_33_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13018_ _05022_ _04516_ _05023_ _05024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_182_3766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_182_3777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15273__A1 _05849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17757_ _00827_ clknet_leaf_49_clk tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14969_ _01744_ channels.sample1\[1\] channels.sample2\[1\] _01758_ _06941_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_16708_ _08445_ _08446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_18_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08490_ _01010_ _01019_ _01020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_17688_ _00758_ clknet_leaf_66_clk tt_um_rejunity_sn76489.tone\[1\].gen.counter\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_162_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16639_ _01715_ _08375_ _08378_ _01717_ _00781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_18_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13587__A1 _04238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13587__B2 _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09111_ channels.accum\[0\]\[22\] _01562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_29_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16525__A1 _08238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09042_ _01491_ _01485_ _01500_ _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_44_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14000__A2 _05954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10573__A1 _02359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15736__I _07636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09944_ channels.freq3\[10\] _02248_ _02243_ _02253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15500__A2 _06910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09734__I _02104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08518__A1 _01024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09875_ _02155_ _02201_ _02204_ _00202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10325__A1 _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08826_ _01298_ _01299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14067__A2 _03377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08757_ _01191_ _01232_ _01237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_169_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13814__A2 _05723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08688_ _01171_ _01172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_75_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15567__A2 _07504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_101_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10650_ _02642_ _02823_ _02908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_81_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09309_ _01730_ _01731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10581_ _02824_ _02840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_180_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09909__I _02226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12320_ _04325_ _04326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_23_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12002__A1 _03925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12251_ _04218_ _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_32_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11202_ filters.sample_filtered\[11\] _03415_ _03416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_121_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12182_ _03183_ _04188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_147_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_147_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11133_ _03345_ _03346_ _03350_ _03229_ _03351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_102_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16990_ _00069_ clknet_leaf_154_clk channels.accum\[0\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_164_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15941_ _07822_ _07823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_11064_ _03285_ _03286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10015_ _02290_ _02302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_125_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15872_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[0\] _07746_ _07754_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_125_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_160_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17611_ _00681_ clknet_leaf_133_clk channels.env_counter\[3\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14823_ _06777_ _06807_ _06808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_99_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13805__A2 _05807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17542_ _00612_ clknet_leaf_243_clk filters.low\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11966_ channels.env_counter\[2\]\[7\] _04030_ _04042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14754_ _06743_ _06744_ _06745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13705_ _05620_ _05621_ _05709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10917_ _03154_ _03104_ _03157_ _00291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_17_Left_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_14685_ _06675_ _06679_ _06680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_17473_ _00543_ clknet_leaf_27_clk filters.band\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__16755__A1 _08449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11897_ _03745_ _03980_ _03981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_16424_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[13\] _08220_ _08229_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_157_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13636_ _05577_ _05640_ _05641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_39_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10848_ _03058_ _03073_ _03100_ _03101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14725__I _06717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13567_ _05503_ _05506_ _05571_ _05572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16355_ channels.ch3_env\[0\] _08179_ _08180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10779_ _03030_ _03032_ _03034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12518_ _03273_ _04243_ _04296_ _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_81_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15306_ _07263_ _07264_ _07265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16286_ _02103_ _07838_ _00676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13498_ filters.high\[20\] filters.band\[20\] _03186_ _05504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_112_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12449_ _04312_ _04449_ _04321_ _04453_ _04455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_15237_ _07176_ _07191_ _07199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15168_ _07125_ _07128_ _07132_ _07133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_22_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14119_ _04801_ _04927_ _06119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_61_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15099_ _07053_ _05421_ _07065_ _07066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__14297__A2 _06285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10307__A1 _01470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09660_ channels.sus_rel2\[6\] _01869_ _02001_ channels.freq2\[6\] _02045_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_94_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14049__A2 _05078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08611_ _01116_ _00022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_136_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09591_ _01874_ _01975_ _01976_ _01978_ _01979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_171_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08542_ _01050_ _01048_ _01055_ _01056_ _00007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_82_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08473_ net7 net16 _01003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__12480__A1 _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13980__A1 _05560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09025_ _01476_ _01474_ _01483_ _01485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_115_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12155__I _04160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16850__I _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08739__A1 _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09087__S1 _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13583__I1 filters.band\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09927_ _01813_ _02240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_102_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_142_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09858_ _02123_ _01830_ _02193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_176_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_142_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08911__A1 _01377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08809_ _01281_ _01282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09789_ channels.sus_rel1\[0\] _02143_ _02138_ _02144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_38_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11820_ _03909_ _03911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13799__A1 _04694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14460__A2 _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output29_I net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11751_ _01166_ _03842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_68_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__16737__A1 _08449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_80_clk clknet_5_9__leaf_clk clknet_leaf_80_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_165_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10702_ _02952_ _02958_ _02959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_14470_ _06458_ _06466_ _06467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_49_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11682_ _03539_ _02711_ _03131_ _03766_ _03772_ _03773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_181_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14212__A2 _05049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13421_ _05405_ _05415_ _05427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_165_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10633_ _02839_ _02868_ _02890_ _02891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_113_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16140_ _08014_ _07961_ _08016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08978__A1 channels.freq2\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08978__B2 channels.freq1\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13352_ _05303_ _05332_ _05357_ _05358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_23_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10564_ _02823_ _02824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10785__A1 _03039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12303_ _04308_ _04309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_16071_ spi_dac_i.spi_dat_buff_1\[2\] _07726_ _07950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_118_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13283_ _05098_ net45 _05288_ _05289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_121_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10495_ _02594_ _02645_ _02756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13318__A4 _04804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09078__S1 _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15022_ _06986_ _06991_ _06992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13723__A1 _05631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12526__A2 _04245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12234_ _03246_ _03193_ _03249_ filters.high\[2\] _04240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_4
XANTENNA__14280__I _06168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12165_ filters.res_lut\[3\] _04170_ _04171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_20_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14279__A2 _06277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11116_ _03210_ _03335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_120_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16973_ _00052_ clknet_leaf_191_clk channels.exp_counter\[2\]\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12096_ _04129_ _00498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15924_ _07783_ _07805_ _07806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_11047_ _03190_ _03193_ _03196_ _03269_ _03270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_36_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput9 bus_in[1] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15855_ _07724_ _07733_ _07738_ _07739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14806_ filters.band\[19\] _06785_ _06763_ _06793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_87_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15786_ _06801_ _07677_ _07688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12998_ _04996_ _05001_ _05003_ _05004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_59_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17525_ _00595_ clknet_leaf_20_clk filters.sample_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__16728__A1 _01806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14737_ _03440_ _06508_ _06729_ _06610_ _00539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_11949_ _03866_ _04023_ _04028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_143_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_177_3665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_71_clk clknet_5_14__leaf_clk clknet_leaf_71_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_59_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_177_3676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_1230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17456_ _00526_ clknet_leaf_0_clk filters.band\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_145_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14668_ _06456_ _06473_ _06663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16407_ _08215_ _08216_ _08211_ _00722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_129_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_138_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13619_ _05487_ _05624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_171_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17387_ _00457_ clknet_leaf_149_clk channels.env_counter\[2\]\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14599_ _06534_ _06594_ _06595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_41_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08969__A1 _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12765__A2 _04766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16338_ _03978_ _08165_ _08169_ _00700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16269_ _08129_ _08131_ _00669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13309__A4 _04803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13714__A1 _05629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09712_ _01819_ _02081_ _02087_ _00156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_87_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09643_ channels.sample3\[9\] _02029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13534__I _04159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09574_ _01933_ _01962_ _00143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_136_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08525_ _01025_ _01050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12453__A1 _03273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_62_clk clknet_5_11__leaf_clk clknet_leaf_62_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_72_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13953__A1 _05950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_98_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09008_ channels.accum\[0\]\[12\] channels.accum\[1\]\[12\] channels.accum\[2\]\[12\]
+ channels.accum\[3\]\[12\] _01140_ _01154_ _01469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10280_ _02382_ _02541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_131_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12613__I _04498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14130__A1 _04371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13970_ _05968_ _05971_ _05972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12921_ _04926_ _04927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12692__A1 _04694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12692__B2 _04697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15640_ _06978_ _07573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14969__B1 channels.sample2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12852_ _04739_ _04858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_69_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11803_ _03893_ _03894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_159_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15571_ _07507_ _07508_ _07509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12783_ _04721_ _04722_ _04789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_84_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11247__A2 _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_53_clk clknet_5_10__leaf_clk clknet_leaf_53_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_56_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17310_ _00380_ clknet_leaf_156_clk channels.accum\[1\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11734_ _03814_ _03824_ _03825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12995__A2 _05000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14522_ _06412_ _06470_ _06518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_138_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_155_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17241_ _00311_ clknet_leaf_11_clk filters.sample_filtered\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11665_ _03530_ _03531_ _03756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14453_ _06448_ _06449_ _06450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_172_3573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13404_ _04876_ _04934_ _05410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_10616_ _02868_ _02874_ _02875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_172_3584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17172_ _00242_ clknet_leaf_125_clk channels.atk_dec3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14384_ _06379_ _06381_ _06382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_92_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11596_ _03666_ _03696_ _03702_ _00425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10758__A1 _01927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12009__B _01032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16123_ _07996_ _07999_ _08000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13335_ _05251_ _05339_ _05340_ _05341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_24_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10547_ _02583_ _02590_ _02807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_45_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16054_ _07767_ _07933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_13266_ _05171_ _05190_ _05272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10478_ _02612_ _02650_ _02739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13619__I _05487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12217_ _03200_ _04216_ _04222_ _04223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_15005_ _06958_ _06975_ _06952_ _06976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13197_ _05199_ _05201_ _05202_ _05203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_clkbuf_leaf_232_clk_I clknet_5_17__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17208__CLK clknet_5_24__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12148_ channels.accum\[3\]\[22\] _04156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10043__I _02293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12079_ _04106_ _04120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16956_ _00035_ clknet_leaf_212_clk channels.lfsr\[3\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15907_ _07786_ _07788_ _07789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_247_clk_I clknet_5_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_179_3705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_139_Right_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16887_ _01196_ _00955_ _00959_ _00964_ _00971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_78_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15838_ spi_dac_i.counter\[3\] _07724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14424__A2 _06027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13227__A3 _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15769_ _03468_ _07670_ _07671_ _07676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_44_clk clknet_5_2__leaf_clk clknet_leaf_44_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_75_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17508_ _00578_ clknet_leaf_247_clk filters.high\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09290_ channels.lfsr\[0\]\[21\] _01717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12986__A2 _04991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15502__C _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14188__A1 _03330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17439_ _00509_ clknet_leaf_169_clk channels.accum\[3\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_172_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_179_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15688__A1 filters.sample_buff\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12910__A2 _04856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_106_Right_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09626_ channels.freq1\[4\] _02011_ _02012_ channels.pw3\[4\] _02013_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_179_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09557_ channels.sus_rel1\[2\] _01899_ _01939_ channels.sample3\[6\] _01945_ _01946_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_78_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08508_ _01031_ _01036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_38_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09488_ _01856_ _01824_ _01853_ _01879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_77_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14179__A1 _03330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11450_ _03607_ _03603_ _01448_ _03604_ _00374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_19_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_110_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10401_ _02561_ _02662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_115_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09150__S0 _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11381_ _02357_ _03566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_132_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_150_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15679__A1 filters.sample_buff\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_150_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13120_ _05122_ _05125_ _05126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10332_ _02592_ _02535_ _02513_ _02593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_131_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13051_ _04629_ _05054_ _05056_ _05057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_111_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10263_ _02508_ _02524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_108_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12002_ _03925_ _04070_ _03935_ _04071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_178_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10194_ _02427_ _02455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_100_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16810_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[3\] _00907_ _00912_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15851__A1 _07721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16741_ _08450_ _00863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13953_ _05950_ _05954_ _05955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09530__A1 channels.ch3_env\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12904_ _04852_ _04857_ _04910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08964__S0 _01148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16672_ _08411_ _08415_ _08281_ _08417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13884_ _05884_ _05885_ _05886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_88_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15623_ _07548_ _07546_ _07556_ _07557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_12835_ _04732_ _04736_ _04841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_115_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_26_clk clknet_5_4__leaf_clk clknet_leaf_26_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_29_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_174_3613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15554_ _07491_ _07492_ _07493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_139_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12766_ _04763_ _04770_ _04771_ _04772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14505_ _06499_ _06501_ _06502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11717_ _03757_ _03806_ _03807_ _03808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_139_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15485_ _06891_ _06719_ _07429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12697_ _04257_ _04703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_83_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17224_ _00294_ clknet_leaf_169_clk channels.sample2\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_11648_ _03738_ _03740_ _00439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14436_ _06339_ _06340_ _06433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_65_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput12 bus_in[4] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_181_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17155_ _00225_ clknet_leaf_141_clk channels.freq3\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09597__B2 channels.pw2\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14590__A1 _05624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11579_ channels.freq3\[5\] _03688_ _03690_ _03692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14367_ _06363_ _06364_ _06365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16106_ _07747_ _07983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13318_ _04695_ _04729_ _05220_ _04804_ _05324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__17030__CLK clknet_5_18__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17086_ _00156_ clknet_leaf_109_clk channels.freq1\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_150_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14298_ _06287_ _06179_ _06293_ _06285_ _06296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA_clkbuf_leaf_171_clk_I clknet_5_24__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14342__A1 _04318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16037_ _07848_ _07863_ _07917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__12253__I _04258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13249_ _05250_ _05254_ _05255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_62_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_51_clk_I clknet_5_10__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08790_ _01250_ _01263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_23_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_186_clk_I clknet_5_22__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14645__A2 _04576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16939_ _00018_ clknet_leaf_220_clk channels.lfsr\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_66_clk_I clknet_5_11__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09521__A1 channels.ctrl_reg2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10131__A2 channels.pw2\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09411_ _01006_ _01805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_133_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_177_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09342_ _01744_ _01745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_177_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12959__A2 _04420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09273_ channels.lfsr\[1\]\[18\] _01703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_30_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_124_clk_I clknet_5_27__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13908__A1 _04406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13908__B2 _04929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09588__A1 channels.freq3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14581__A1 _04802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12187__A3 _04192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_95_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer20_I _05151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09737__I _02106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_139_clk_I clknet_5_31__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_19_clk_I clknet_5_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12895__A1 _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08988_ _01442_ _01443_ _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16881__I0 _00966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12647__A1 _04535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10950_ channels.sample1\[10\] _01261_ _03177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_27_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09609_ _01847_ _01996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10881_ _03131_ _02940_ _03132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12620_ _04623_ _04624_ _04626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__09276__B1 _01705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12551_ _04362_ _04428_ _04309_ _04557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_81_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_152_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11502_ _02326_ _03632_ _03637_ _00396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_53_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12482_ _03238_ _03182_ _04188_ _03410_ _04488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_15270_ _07227_ _07230_ _07231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_108_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09579__A1 filters.res_filt\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14572__A1 _04326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14221_ _06116_ _06117_ _06220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_11433_ channels.accum\[1\]\[4\] _03597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09579__B2 channels.freq2\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14152_ _04258_ _05504_ _06152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_130_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11364_ _01088_ _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13127__A2 _05114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10315_ _02575_ _02576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13103_ _05104_ _05105_ _05108_ _05109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_21_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14083_ _06000_ _06057_ _06083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_11295_ _03499_ _03500_ _03501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13034_ _05032_ _05034_ _05040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10246_ _02484_ _02498_ _02386_ _02507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_28_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_167_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09751__A1 channels.ctrl_reg1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10177_ _02434_ _02435_ _02436_ _02437_ _01527_ _02438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__09382__I _01780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15824__A1 _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_128_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17773_ _00843_ clknet_leaf_203_clk channels.exp_periods\[1\]\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14985_ filters.high\[3\] _06955_ _06956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09503__A1 channels.pw1\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09503__B2 channels.freq2\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16724_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[8\] _08454_ _08451_ _08458_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13936_ _04446_ _04766_ _05724_ _05938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_156_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10113__A2 channels.ring_outs\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16655_ _08395_ _08402_ _08403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_158_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13867_ _05864_ _05867_ _05868_ _05869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_69_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15606_ channels.sample2\[7\] _03395_ _07540_ _03232_ _07541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_29_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12818_ _04780_ _04824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16586_ _08358_ _08361_ _08362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13798_ _05512_ _05091_ _05079_ _05800_ _05801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_173_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15537_ channels.sample1\[2\] _03335_ _07477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12749_ _04741_ _04743_ _04755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__12810__A1 filters.cutoff_lut\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15468_ filters.high\[28\] _07030_ _07356_ _07414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_167_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17207_ _00277_ clknet_leaf_173_clk channels.sample3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_128_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10991__I _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14419_ _06319_ _06324_ _06416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_114_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15399_ _07342_ _07345_ _07349_ _07350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_170_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17138_ _00208_ clknet_leaf_124_clk channels.atk_dec2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_163_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09990__A1 channels.ctrl_reg3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09960_ _02242_ _02257_ _02263_ _00228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17069_ _00139_ clknet_leaf_98_clk filters.hp vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__16855__A3 _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_6_clk clknet_5_5__leaf_clk clknet_leaf_6_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_100_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_90_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08911_ _01377_ _01378_ _01379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09891_ _01776_ _02215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12877__A1 _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09742__A1 _02110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08842_ _01303_ _01314_ _01315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_100_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12629__A1 _03256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08773_ _01247_ _00053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_174_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11301__A1 _02316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10104__A2 _01230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13841__A3 _05843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13542__I _05546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09325_ _01689_ _01734_ _01735_ _01692_ _00117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12801__A1 _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12158__I _04163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09256_ _01682_ _01683_ _01689_ _01674_ _00094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_173_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_32_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09187_ channels.lfsr\[1\]\[5\] _01630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_172_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09981__A1 channels.ctrl_reg3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13109__A2 _05114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14306__A1 _05877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15503__B1 _03476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10100_ _01282_ _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_11080_ _03300_ _03301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_179_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15418__B _07356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13717__I _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10031_ _02308_ _02310_ _02313_ _00249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09416__B _01809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15806__A1 _07373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14609__A2 _06501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_26__f_clk clknet_3_6_0_clk clknet_5_26__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_145_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15282__A2 _07033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14770_ _04159_ _06760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11982_ _04053_ _04054_ _04055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_106_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09930__I _01818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13721_ _05720_ _05724_ _05725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10933_ channels.sample1\[3\] _03164_ _03167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_123_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_123_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16440_ _08240_ _08241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_168_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13045__A1 _04928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13652_ _05553_ _05642_ _05656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10864_ _03112_ _03115_ _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_151_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12603_ _04563_ _04572_ _04609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_66_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12068__I _04103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16763__I _02101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16371_ channels.ch3_env\[7\] _08185_ _08189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10795_ _02983_ _03010_ _03008_ _03050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13583_ filters.high\[21\] filters.band\[21\] _05179_ _05588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_112_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_171_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15322_ _07278_ _07279_ _07280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_164_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12534_ _04537_ _04165_ _04538_ _04539_ _04540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_82_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15379__I _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15253_ _07211_ _07214_ _07215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12465_ _04470_ _04471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11700__I _03532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09377__I _01776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14204_ _06112_ _06113_ _06203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11416_ channels.accum\[2\]\[21\] _03556_ _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_169_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12396_ _03190_ _03312_ _03196_ filters.high\[10\] _04402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
X_15184_ _07113_ _07117_ _07135_ _07138_ _07148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_111_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10031__A1 _02308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14135_ _06122_ _06134_ _06135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_11347_ _03539_ _03540_ _03541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11278_ _02308_ _03484_ _03486_ _00323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12859__A1 _04200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14066_ _06066_ _06067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_39_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09724__A1 _01767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13017_ _04381_ _04439_ _04496_ _05023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_10229_ _01510_ _02473_ _02490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_182_3756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_5_14__f_clk_I clknet_3_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17756_ _00826_ clknet_leaf_49_clk tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14968_ _01758_ _01744_ channels.sample1\[1\] channels.sample2\[1\] _06940_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__09840__I _02104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16707_ _08441_ _08442_ _08444_ _08445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_18_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13919_ _05836_ _05837_ _05921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_17687_ _00757_ clknet_leaf_66_clk tt_um_rejunity_sn76489.tone\[1\].gen.counter\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_18_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14899_ _06875_ _03476_ _06876_ _06877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16222__A1 _07726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16638_ _01710_ _08375_ _08378_ _01712_ _00780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_29_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16569_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[4\] _08328_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[4\]
+ _08348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_29_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_174_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09110_ _01540_ _01559_ _01561_ _00076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10270__A1 _01305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09041_ _01499_ _01500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12706__I _04711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11610__I _03711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_111_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10022__A1 _02240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10573__A2 _02831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09943_ _02187_ _02252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_1_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12441__I _04446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13511__A2 _05516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09874_ channels.ctrl_reg2\[5\] _02202_ _02199_ _02204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10325__A2 _02377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08825_ _01270_ _01297_ _01298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_174_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15752__I _07663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16461__A1 _08136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08756_ _01236_ _00047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input10_I bus_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09750__I _02106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08687_ _01170_ _01171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_138_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_101_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11589__A1 channels.pw3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09308_ _01725_ _01730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10580_ _02703_ _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_81_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10261__A1 _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09239_ _01669_ _01659_ _01673_ _01674_ _00092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_35_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11520__I _03641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12250_ _03254_ _04226_ _04255_ _04256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_107_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10013__A1 _02299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11201_ _03410_ _03233_ _03414_ _03415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_31_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12181_ _04186_ _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13750__A2 _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_147_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11132_ _03349_ _03350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_147_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_164_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_164_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15940_ _07821_ _07818_ _07822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11063_ _03246_ _03283_ _03249_ _03284_ _03285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XANTENNA__10316__A2 _02569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11513__A1 channels.pw1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10014_ _02290_ _02301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15871_ _07749_ _07751_ _07752_ _07753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_125_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17610_ _00680_ clknet_leaf_133_clk channels.env_counter\[3\]\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15255__A2 _07216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14822_ filters.low\[21\] filters.band\[21\] _06073_ _06807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_99_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17541_ _00611_ clknet_leaf_5_clk filters.low\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14753_ _06732_ _06736_ _06744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11965_ _03935_ _04039_ _04040_ _04041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_25_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_129_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13704_ _05611_ _05706_ _05707_ _05708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_169_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17472_ _00542_ clknet_leaf_245_clk filters.band\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10916_ channels.sample2\[8\] _03156_ _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14684_ _06676_ _06677_ _06678_ _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_168_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11896_ _03754_ _03543_ _03946_ _03980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_128_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16423_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[12\] _08223_ _08228_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13635_ _05579_ _05639_ _05640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_67_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_156_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10847_ _03061_ _03072_ _03100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16354_ _08178_ _08179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_171_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13566_ _04597_ _05570_ _05507_ _05571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_87_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10778_ _03030_ _03032_ _03033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_82_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15305_ _07260_ _07262_ _07264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_125_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12517_ _03333_ _04293_ _04522_ _04523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_16285_ _08140_ _08141_ _07740_ _00675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13497_ _04295_ _05279_ _05503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_164_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15236_ _07164_ _07168_ _07198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_180_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12448_ _04449_ _04322_ _04453_ _04312_ _04454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_152_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_75_Right_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09945__A1 _02252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10046__I _02154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15167_ _07129_ _07130_ _07131_ _07132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_10_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12379_ _04384_ _04385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_14118_ _06116_ _06117_ _06118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_1_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15098_ _05417_ _05420_ _07065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_120_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14049_ _04372_ _05078_ _06050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input2_I addr[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11504__A1 _02328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_158_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_230_clk clknet_5_17__leaf_clk clknet_leaf_230_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_2_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08610_ channels.lfsr\[3\]\[9\] _01116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09590_ channels.ctrl_reg1\[3\] _01941_ _01903_ _01977_ _01978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_59_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_84_Right_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17739_ _00809_ clknet_leaf_53_clk tt_um_rejunity_sn76489.control_tone_freq\[0\]\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08541_ _01040_ _01050_ _01045_ _00006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08472_ _01000_ _01001_ _01002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_175_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_46_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09024_ _01476_ _01474_ _01483_ _01484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_116_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_93_Right_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_170_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09926_ _02238_ _02235_ _02239_ _00218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13496__A1 _04525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09857_ _02191_ _02181_ _02192_ _02103_ _00196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_142_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_221_clk clknet_5_21__leaf_clk clknet_leaf_221_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08808_ _01280_ _01281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XPHY_EDGE_ROW_0_Left_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09788_ _02141_ _02143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08739_ _01169_ _01206_ _01222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_120_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11750_ _03836_ _03840_ _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_83_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10701_ _02953_ _02957_ _02958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_55_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11681_ _03768_ _03088_ _03771_ _03747_ _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_138_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13420_ _05378_ _05404_ _05426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_153_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10632_ _02873_ _02890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_157_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13351_ _05335_ _05356_ _05357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_10563_ _02768_ _02820_ _02822_ _02774_ _02823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_52_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12302_ _04213_ _04306_ _04307_ _04308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16070_ _07926_ _07947_ _07721_ _07949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_118_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13282_ _05196_ _05286_ _05288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10494_ _02641_ _02501_ _02755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15021_ _06989_ _06990_ _06991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__13723__A2 _05632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12233_ _03200_ _04216_ _04238_ _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_20_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12164_ _04169_ _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_9_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13177__I _04858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11115_ _03329_ _03218_ _03333_ _03228_ _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_16972_ _00051_ clknet_5_23__leaf_clk channels.exp_counter\[2\]\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12095_ _03545_ channels.adsr_state\[2\]\[0\] _04128_ _04129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15923_ _07789_ _07796_ _07804_ _07805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11046_ filters.band\[2\] _03269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
Xclkbuf_leaf_212_clk clknet_5_20__leaf_clk clknet_leaf_212_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_21_1298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15854_ spi_dac_i.counter\[4\] _07733_ _07724_ _07738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13239__A1 _05157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14805_ _06748_ _06791_ _06792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_15785_ _07686_ _07687_ _00629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_153_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12997_ _05002_ _05000_ _05003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17524_ _00594_ clknet_leaf_19_clk filters.sample_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14736_ _06403_ _06728_ _06729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11948_ _04006_ _04027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_177_3666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_177_3677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17455_ _00525_ clknet_leaf_188_clk channels.accum\[3\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14667_ _06655_ _06658_ _06661_ _06662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_157_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11879_ channels.env_vol\[0\]\[4\] _03965_ _03966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16406_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[8\] _08209_ _08216_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_138_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13618_ _05619_ _05622_ _05623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_171_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17386_ _00456_ clknet_leaf_136_clk channels.env_counter\[2\]\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_138_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14598_ _06537_ _06593_ _06594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_89_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16337_ channels.env_vol\[1\]\[6\] _08166_ _08169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13549_ _05444_ _05454_ _05554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_41_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09091__A1 _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16268_ filters.sample_buff\[10\] _08125_ _08130_ spi_dac_i.spi_dat_buff_0\[6\] spi_dac_i.spi_dat_buff_0\[7\]
+ _08127_ _08131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_113_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_164_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09918__A1 _02215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15219_ _07181_ _07182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_164_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16199_ _08057_ _08072_ _08073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_61_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12920__S _03185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09711_ channels.freq1\[15\] _02082_ _02084_ _02087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_87_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_203_clk clknet_5_21__leaf_clk clknet_leaf_203_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09642_ _02024_ _02025_ _02026_ _02027_ _02028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_179_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09573_ _01934_ net24 _01947_ _01961_ _01962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_117_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08524_ _01049_ _00002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13650__A1 _05527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12453__A2 _04372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13402__A1 _04938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13253__I1 filters.band\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13953__A2 _05954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_36_Left_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09007_ _01466_ _01467_ _01468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_170_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13705__A2 _05621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11716__A1 channels.atk_dec3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11716__B2 channels.atk_dec2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11192__A2 _03385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09909_ _02226_ _02228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14130__A2 _05185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_45_Left_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12920_ filters.high\[15\] filters.band\[15\] _03185_ _04926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__16101__I _07956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08896__A1 channels.freq3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12692__A2 _04281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12851_ _04853_ _04855_ _04856_ _04857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_68_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11802_ _03884_ _03885_ _03887_ _03891_ _03892_ _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_TAPCELL_ROW_159_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15570_ _07499_ _07496_ _07506_ _07508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_159_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12782_ _04721_ _04722_ _04788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_96_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14521_ _06476_ _06487_ _06516_ _06517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11733_ _03823_ _03824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13460__I _04805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17240_ _00310_ clknet_5_7__leaf_clk filters.sample_filtered\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_181_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14452_ _06358_ _06367_ _06449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11664_ _03745_ _03754_ _03755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_25_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_54_Left_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_154_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13403_ _05407_ _05408_ _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_36_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17171_ _00241_ clknet_leaf_125_clk channels.atk_dec3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10615_ _02504_ _02873_ _02874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_172_3574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14383_ _06380_ _04632_ _06381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_172_3585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11595_ channels.pw3\[3\] _03697_ _03698_ _03702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16122_ _07997_ _07998_ _07999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13334_ _04254_ _04470_ _04490_ _04712_ _05340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_3_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10546_ _02750_ _02805_ _02806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__16343__B1 _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16053_ _07777_ _07890_ _07932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13265_ _05087_ _05269_ _05270_ _05271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10477_ _02616_ _02617_ _02737_ _02738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__09385__I net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15004_ _06971_ _06974_ _06975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_12216_ _04221_ _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_13196_ _05138_ _05152_ _05202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16646__A1 _08267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12147_ _04155_ _00523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_63_Left_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10930__A2 _02831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12078_ _04103_ _04119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16955_ _00034_ clknet_leaf_224_clk channels.lfsr\[3\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15906_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[1\] _07787_ _07788_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_159_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11029_ _03252_ _03253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16886_ _01202_ _00938_ _00970_ _00840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_154_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_179_3706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15837_ _07719_ _07723_ _07573_ _00645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_91_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15621__A2 _07554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15768_ _06746_ _07664_ _07675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_17507_ _00577_ clknet_leaf_247_clk filters.high\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14719_ _06689_ _06712_ _06713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_59_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15699_ _07624_ _00606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_72_Left_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_145_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_60_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17438_ _00508_ clknet_leaf_181_clk channels.accum\[3\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_133_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17369_ _00439_ clknet_leaf_165_clk channels.clk_div\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12738__A3 _04743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_141_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_58_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_81_Left_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__16637__A1 _01705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_7__f_clk clknet_3_1_0_clk clknet_5_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10921__A2 _03136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09119__A2 _01566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13871__A1 _05743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09625_ _01896_ _02012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09556_ _01940_ _01942_ _01944_ _01945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_66_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_90_Left_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08507_ _01030_ _01034_ _01035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09487_ channels.ch3_env\[0\] _01877_ _01878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14179__A2 _06177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10400_ _02654_ _02659_ _02660_ _02661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09150__S1 _01154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11380_ _03565_ _03557_ _01395_ _03558_ _00346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_115_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_150_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10331_ _02507_ _02592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10262_ _02509_ _02514_ _02522_ _02523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_13050_ _05052_ _05055_ _05056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__13154__A3 _04375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11796__S0 _03886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12001_ _03920_ _04066_ _04070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__16628__A1 _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10193_ channels.pw2\[2\] _02454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_1296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16740_ _08453_ _08464_ _00862_ _00802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13952_ _05951_ _05952_ _05953_ _05954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__08869__A1 channels.freq2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08869__B2 channels.freq1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13862__A1 _05852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12903_ _04866_ _04909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_16671_ _08411_ _08415_ _08416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__16766__I _03494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13883_ _05440_ _05766_ _05779_ _05885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08964__S1 _01163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15622_ _07555_ _07556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_159_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12834_ _04815_ _04839_ _04840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_119_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13614__A1 _04864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_174_3614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15553_ channels.sample1\[3\] _03400_ _07492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12765_ _04765_ _04766_ _04769_ _04771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_56_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14504_ _03380_ _03378_ _06500_ _06501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_11716_ channels.atk_dec3\[2\] _03782_ _01278_ channels.atk_dec2\[2\] _03785_ _03807_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_12_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15484_ _07427_ _07428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__15367__B2 _07277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12696_ _04388_ _04480_ _04702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17223_ _00293_ clknet_leaf_93_clk channels.sample2\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14435_ _06417_ _06431_ _06432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11647_ _02272_ _03739_ _03740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09046__A1 _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_182_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput13 bus_in[5] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_140_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11928__A1 _01581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17154_ _00224_ clknet_leaf_141_clk channels.freq3\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14366_ _04222_ _05793_ _06364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11578_ _03668_ _03687_ _03691_ _00418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_16105_ _07749_ _07751_ _07982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13317_ _05236_ _05237_ _05322_ _05323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_17085_ _00155_ clknet_leaf_109_clk channels.freq1\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10529_ _02741_ _02780_ _02789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_40_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_172_Right_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14297_ _06294_ _06285_ _06295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_123_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16036_ _07915_ _07916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13248_ _05251_ _05252_ _05253_ _05254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_58_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12353__A1 _04356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13179_ filters.high\[17\] filters.band\[17\] _03186_ _05185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_36_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10903__A2 _02932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10989__I _03204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_53_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16938_ _00017_ clknet_leaf_220_clk channels.lfsr\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13853__A1 _05852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09521__A2 _01830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16869_ _00940_ _00952_ _00956_ _01183_ _00957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_09410_ _01801_ _01802_ _01804_ _00137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10419__A1 _02607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08707__S1 _01172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09341_ filters.filt_1 _01744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13081__A2 _05049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09272_ channels.lfsr\[0\]\[18\] _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13908__A2 _05909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12592__A1 _04468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08796__B1 channels.ctrl_reg1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12444__I _04375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12344__A1 _04252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_73_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14097__A1 _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08987_ _01299_ _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_119_Left_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09608_ channels.ctrl_reg2\[4\] _01974_ _01966_ channels.atk_dec2\[4\] _01994_ _01995_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_108_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10880_ _03088_ _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_35_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09539_ _01924_ _01925_ _01926_ _01928_ _01929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_78_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09276__B2 _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_231_clk_I clknet_5_20__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12550_ _04548_ _04554_ _04555_ _04556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_93_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_152_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16535__B _08318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11501_ channels.freq1\[6\] _03633_ _03634_ _03637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12481_ _04185_ _04487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_47_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14220_ _06217_ _06131_ _06218_ _06219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09579__A2 _01844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11432_ _03160_ _01359_ _03596_ _00367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_128_Left_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08832__I _01142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14572__A2 _05891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_246_clk_I clknet_5_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12583__A1 _04583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16849__A1 _01581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14151_ _05069_ _05350_ _06151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_130_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11363_ _03555_ _00339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13102_ _03199_ _04215_ _05107_ _05108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_10314_ _01687_ _02572_ _02574_ _02575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_14082_ _05984_ _05996_ _06081_ _06082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_104_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11294_ _03497_ _03500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_131_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11138__A2 _03337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13033_ _05029_ _05038_ _05017_ _05039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10245_ _02502_ _02505_ _02506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_167_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10897__A1 channels.sample2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10176_ _02428_ channels.pw2\[5\] _01097_ _02437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__14088__A1 _05440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15824__A2 _04158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_137_Left_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_128_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17772_ _00842_ clknet_leaf_200_clk channels.exp_periods\[1\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14984_ _06952_ _06955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_92_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09503__A2 _01891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16723_ _08456_ _08446_ _08457_ _00797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13935_ _05799_ _05808_ _05936_ _05937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_16654_ _08397_ _08401_ _08402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_158_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13866_ _05852_ _05855_ _05868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15605_ _03358_ _07538_ _07539_ _06710_ _07540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_12817_ _03271_ _04242_ _04784_ _04823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_16585_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[7\] _08329_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[7\]
+ _08361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13797_ _04471_ _05800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15536_ channels.sample2\[2\] _03346_ _07475_ _03229_ _07476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_12748_ _04286_ _04753_ _04754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10049__I _01813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15467_ _07408_ _07412_ _07413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_5_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14012__A1 _04694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12679_ _04551_ _04553_ _04548_ _04685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__08490__A2 _01019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17206_ _00276_ clknet_leaf_174_clk channels.sample3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14418_ _06413_ _06414_ _06415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15398_ _07348_ _07344_ _07349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17137_ _00207_ clknet_leaf_127_clk channels.atk_dec2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14349_ _06314_ _06346_ _06347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_123_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_38_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17068_ _00138_ clknet_leaf_99_clk filters.bp vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__13118__A3 _04450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15512__A1 channels.sample3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16019_ _07897_ _07898_ _07899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08910_ channels.accum\[0\]\[5\] channels.accum\[1\]\[5\] channels.accum\[2\]\[5\]
+ channels.accum\[3\]\[5\] _01147_ _01161_ _01378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_90_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09890_ _02188_ _02210_ _02214_ _00207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_85_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12877__A2 _04215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08841_ _01304_ _01310_ _01313_ _01314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14079__A1 _03314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11608__I _01740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15815__A2 _07697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08772_ channels.exp_counter\[2\]\[4\] _01245_ _01238_ _01084_ _01247_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12629__A2 _04566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09050__S0 _00009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15579__A1 channels.sample2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12439__I _04444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14251__A1 _06236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09324_ _01681_ _01734_ _01735_ _01685_ _00116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_146_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12801__A2 _04802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09255_ _01684_ _01685_ _01675_ _01686_ _01144_ _01688_ _01689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_111_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14929__I1 filters.band\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08481__A2 _01003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09186_ channels.lfsr\[0\]\[5\] _01629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_69_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_181_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12565__A1 _04297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15503__A1 _01748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15503__B2 _01762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_179_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10030_ channels.sus_rel3\[0\] _02311_ _02312_ _02313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_179_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10879__A1 _03128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13817__A1 _05158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11981_ _03914_ _03843_ _04039_ _04054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09497__A1 channels.pw1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09497__B2 channels.freq1\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13720_ _05722_ _05723_ _05724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_169_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10932_ _03162_ _02880_ _03166_ _00297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_123_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13651_ _05553_ _05642_ _05655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_170_clk_I clknet_5_24__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10863_ _03113_ _03114_ _03115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12602_ _04595_ _04606_ _04607_ _04608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_16370_ _03978_ _08184_ _08188_ _00713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_50_clk_I clknet_5_10__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13582_ _04294_ _05186_ _05587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10794_ _03047_ _03048_ _03049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_66_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15321_ filters.low\[16\] _06176_ _07279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_93_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12533_ _04523_ _04524_ _04539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_109_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_185_clk_I clknet_5_22__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15252_ _07212_ _07213_ _07214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12464_ _04257_ _04470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_87_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14203_ _06110_ _06111_ _06202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11415_ _03586_ _03581_ _01552_ _03582_ _00360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_34_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15183_ _07135_ _07138_ _07147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_169_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12395_ _04400_ _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_169_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14134_ _06125_ _06133_ _06134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11346_ _03028_ _03540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_132_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13505__B1 _04946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10582__A3 _02840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14065_ _03375_ _06066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_11277_ filters.cutoff_lut\[6\] _03484_ _03485_ _03486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12859__A2 _04864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13016_ _04381_ _04439_ _04496_ _05022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10228_ _02463_ _02488_ _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_182_3757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_123_clk_I clknet_5_30__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10159_ _02410_ _02411_ _02412_ _02420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__16470__A2 _08263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15273__A3 _07233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17755_ _00825_ clknet_leaf_49_clk tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14967_ _04520_ _04692_ _06939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_16706_ _08443_ _01816_ _03494_ _08444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__11295__A1 _03499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10098__A2 _01245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13918_ _05832_ _05840_ _05919_ _05920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_17686_ _00756_ clknet_leaf_66_clk tt_um_rejunity_sn76489.tone\[1\].gen.counter\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14898_ _06614_ _03475_ _06876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_18_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_138_clk_I clknet_5_31__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16637_ _01705_ _08388_ _08389_ _01707_ _00779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_71_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13849_ _05849_ _05851_ _05852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_76_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_18_clk_I clknet_5_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16568_ _08243_ _08347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_128_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15519_ _07382_ _07460_ _00590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_17_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16499_ _08243_ _08289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09660__A1 channels.sus_rel2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09040_ _01494_ _01498_ _01499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_127_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_5_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11112__B _03330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09942_ _02250_ _02247_ _02251_ _00222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_110_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09873_ _02150_ _02201_ _02203_ _00201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08824_ _01271_ _01283_ _01296_ _01297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08755_ channels.exp_counter\[1\]\[3\] _01230_ _01235_ _01220_ _01236_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10089__A2 _02351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_68_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08686_ _01165_ _01170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_136_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_68_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14224__A1 _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_101_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09100__B1 _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09307_ _01728_ _01729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12786__A1 _04311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_81_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12250__A3 _04255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09238_ _01626_ _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09403__A1 filters.mode_vol\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09169_ _01612_ _01613_ _01600_ _01614_ _01141_ _01155_ _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_47_1230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11200_ _03411_ _03223_ _03413_ _03233_ _03414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_181_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12180_ _04185_ _04186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_31_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13728__I _05731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_147_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11131_ _03348_ _03349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_147_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11062_ filters.band\[3\] _03284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_10013_ _02299_ _02291_ _02300_ _00244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_15870_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[0\] _07749_ _07752_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_125_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_5_6__f_clk_I clknet_3_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14821_ _06769_ _06794_ _06805_ _06806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_1273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13463__I _04737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11277__A1 filters.cutoff_lut\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17540_ _00610_ clknet_leaf_5_clk filters.low\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14752_ _06722_ _06731_ _06743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11964_ _03854_ _04032_ _03903_ _04040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_153_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13703_ _05612_ _05613_ _05707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__12079__I _04106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10915_ _03149_ _03156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17471_ _00541_ clknet_leaf_21_clk filters.band\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14683_ _06441_ _06676_ _06677_ _06678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_157_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11895_ _03960_ _03978_ _03979_ _00447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14215__A1 _06211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16422_ _08226_ _08227_ _08222_ _00726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_157_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13634_ _05602_ _05638_ _05639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10846_ _03094_ _03098_ _03099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_6_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12777__A1 filters.cutoff_lut\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16353_ _02356_ _03936_ _01821_ _08178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13565_ _05501_ _05570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_27_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10777_ _03031_ _02777_ _03032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09388__I net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15304_ _07260_ _07262_ _07263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_124_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12516_ net60 _04522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16284_ spi_dac_i.spi_dat_buff_0\[11\] _08117_ _08141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13496_ _04525_ _05501_ _05502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15235_ _07146_ _07149_ _07196_ _07169_ _07197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_12447_ _04452_ _04453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_140_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11201__A1 _03410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15166_ _01747_ channels.sample1\[8\] _07131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12378_ _04162_ _03315_ _04384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_0_1_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14117_ _04803_ _04861_ _06117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11329_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[1\] _03523_ _03517_ _03526_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15097_ _06913_ _07064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_157_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14048_ _04377_ _05074_ _06049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09851__I _02187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10997__I _03221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15999_ _07747_ _07878_ _07879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08540_ _01060_ _00005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17738_ _00808_ clknet_leaf_53_clk tt_um_rejunity_sn76489.control_tone_freq\[0\]\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08467__I net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08471_ net2 net1 _01001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17669_ _00739_ clknet_leaf_80_clk tt_um_rejunity_sn76489.tone\[2\].gen.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14206__A1 _04750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_46_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_63_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09633__A1 filters.cutoff_lut\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11621__I _03711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09298__I _01032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13041__C _04993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09023_ _01479_ _01482_ _01483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_26_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13193__A1 _05138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09925_ channels.sus_rel2\[5\] _02236_ _02232_ _02239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09856_ _02098_ _02182_ _02192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_176_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08807_ _01279_ _01280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09787_ _02141_ _02142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11259__A1 _03468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08738_ _01221_ _00044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_120_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15712__B _07356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08669_ _00010_ _01153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09872__A1 channels.ctrl_reg2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10700_ _02954_ _02956_ _02957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_178_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11680_ _03769_ _03770_ _03771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_37_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10631_ _02687_ _02840_ _02866_ _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_48_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12627__I _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10234__A2 channels.ctrl_reg2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13350_ _05338_ _05355_ _05356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_148_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10562_ _01556_ _02770_ _02821_ _02822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_91_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16543__B _08313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12301_ _04249_ _04284_ _04305_ _04307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_84_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13281_ _05196_ _05286_ _05287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_101_Left_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_118_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10493_ _02748_ _02749_ _02753_ _02754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__16370__A1 _03978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15020_ _01768_ channels.sample3\[3\] _06990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12232_ _04237_ _04238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_31_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14063__B net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12931__A1 _04644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12163_ _04168_ _04169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_9_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11114_ _03332_ _03333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_102_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16971_ _00050_ clknet_leaf_194_clk channels.exp_counter\[2\]\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12094_ _01240_ _03551_ _01931_ _04128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_15922_ _07803_ _07804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11498__A1 _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11045_ filters.low\[2\] _03268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_21_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15853_ _07737_ _00647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_110_Left_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10170__A1 channels.pw1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14804_ _06788_ _06790_ _06791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12996_ _04998_ _05002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_15784_ filters.low\[19\] _07682_ _07684_ _07687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12998__A1 _04996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17523_ _00593_ clknet_leaf_20_clk filters.sample_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11947_ _04008_ _04025_ _04026_ _00452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14735_ _06724_ _06727_ _06728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09863__A1 channels.ctrl_reg2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_177_3667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14666_ _06534_ _06659_ _06660_ _06661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_17454_ _00524_ clknet_leaf_155_clk channels.accum\[3\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11878_ _03941_ _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16405_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[7\] _08212_ _08215_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13617_ _05620_ _05621_ _05622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_131_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10829_ _03077_ _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_17385_ _00455_ clknet_5_31__leaf_clk channels.env_counter\[2\]\[6\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_138_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09615__A1 channels.sus_rel2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14597_ _06560_ _06592_ _06593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13548_ _05435_ _05551_ _05552_ _05553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_41_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16336_ _03974_ _08165_ _08168_ _00699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10057__I _02330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16267_ _08116_ _08130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_140_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13479_ _04477_ _04884_ _05485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16361__A1 channels.ch3_env\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15164__A2 channels.sample3\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09846__I _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15218_ _07158_ _07159_ _07180_ _07181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16198_ _08069_ _08071_ _08072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_26_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12922__A1 _04487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15149_ _03345_ _07077_ _07115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_77_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14675__A1 _05268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09710_ _01814_ _02081_ _02086_ _00155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11489__A1 _03511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09641_ channels.pw1\[5\] _02003_ _02004_ channels.ctrl_reg1\[5\] _02027_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_136_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09572_ _01875_ _01949_ _01953_ _01960_ _01961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_93_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14978__A2 _06949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08523_ _01047_ _00132_ _01048_ _01049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13650__A2 _05530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12447__I _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_175_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11413__A1 _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09006_ channels.freq2\[12\] _01279_ _01292_ channels.freq1\[12\] _01467_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09908_ _02226_ _02227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09491__I _01881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09839_ _02160_ _02170_ _02178_ _00192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12850_ _03349_ net68 _04192_ _04856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__14969__A2 channels.sample1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11801_ channels.env_counter\[0\]\[10\] channels.env_counter\[1\]\[10\] channels.env_counter\[2\]\[10\]
+ channels.env_counter\[3\]\[10\] _03886_ _01170_ _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_96_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12781_ _04778_ _04786_ _04787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09845__A1 _02179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_159_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14520_ _06479_ _06486_ _06516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11732_ _03819_ _03821_ _03822_ _03533_ _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_56_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08835__I _01307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14451_ _06361_ _06366_ _06448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11663_ _03535_ _03751_ _03753_ _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_181_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_154_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_153_Right_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_138_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11261__I _03470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13402_ _04938_ _04949_ _05408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17170_ _00240_ clknet_leaf_144_clk channels.ctrl_reg3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10614_ _02872_ _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_107_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14382_ filters.band\[26\] _06380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_172_3575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11594_ _03664_ _03696_ _03701_ _00424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_24_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09073__A2 _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16121_ _07963_ _07967_ _07998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13333_ net68 _04490_ _04712_ _04703_ _05339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10545_ _02529_ _02573_ _02804_ _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xclkbuf_leaf_130_clk clknet_5_30__leaf_clk clknet_leaf_130_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_51_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16052_ _07784_ _07930_ _07885_ _07887_ _07883_ _07931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_106_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13264_ _04765_ _05268_ _05090_ _05270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_33_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08570__I _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10476_ _02703_ _02618_ _02624_ _02737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_121_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12904__A1 _04852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15003_ _06948_ _06972_ _06973_ _06974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_12215_ _04220_ _04221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_32_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13195_ _05200_ _05157_ _05163_ _05201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_20_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12146_ channels.accum\[3\]\[21\] _04155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12077_ _04041_ _04113_ _04118_ _00490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16954_ _00033_ clknet_leaf_232_clk channels.lfsr\[3\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15905_ tt_um_rejunity_sn76489.chan\[0\].attenuation.in _07787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_11028_ _03247_ _03248_ _03250_ _03251_ _03252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_95_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16885_ _00939_ _00969_ _00970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_197_clk clknet_5_23__leaf_clk clknet_leaf_197_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_179_3707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15836_ _07720_ _04776_ _07722_ _07723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__16448__B _08098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09836__A1 channels.freq2\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12979_ _04978_ _04979_ _04985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_15767_ _07673_ _07674_ _00624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_129_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17506_ _00576_ clknet_leaf_248_clk filters.high\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11643__A1 _03728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14718_ _03423_ _06710_ _06711_ _06712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_15698_ channels.exp_periods\[3\]\[1\] _07624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_87_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_60_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17437_ _00507_ clknet_leaf_180_clk channels.accum\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14649_ _06551_ _06556_ _06644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_60_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_120_Right_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_157_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17368_ _00438_ clknet_leaf_85_clk channels.clk_div\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_27_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16319_ _02363_ _03937_ _08157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_121_clk clknet_5_27__leaf_clk clknet_leaf_121_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_15_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16334__A1 _03964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17299_ _00369_ clknet_leaf_179_clk channels.accum\[1\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13148__A1 _05122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08480__I net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_58_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10382__A1 _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14648__A1 _05509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13320__A1 _04323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_188_clk clknet_5_19__leaf_clk clknet_leaf_188_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_173_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13871__A2 _05746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09624_ _01954_ _02011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11882__A1 _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09555_ filters.cutoff_lut\[8\] _01849_ _01943_ channels.sus_rel3\[2\] _01944_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08506_ _01031_ _01033_ _01034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09486_ _01876_ _01877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08655__I _01138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_22_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16573__A1 _08314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_92_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17747__CLK clknet_5_8__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_112_clk clknet_5_15__leaf_clk clknet_leaf_112_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_144_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_150_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10330_ _02522_ _02590_ _02591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10261_ _01688_ _02517_ _02521_ _02522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_12000_ _04007_ _04068_ _04069_ _00462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08566__A1 _01070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12362__A2 _03270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11796__S1 _01166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10192_ _01541_ _02433_ _02443_ _02451_ _02452_ _01533_ _02453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
XANTENNA__09515__B1 _01905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13951_ _04392_ _05347_ _05953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_179_clk clknet_5_18__leaf_clk clknet_leaf_179_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12902_ _04852_ _04857_ _04908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16670_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[4\] _08399_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[4\]
+ _08415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13882_ _04667_ _05883_ _05777_ _05884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10676__A2 _02932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15621_ filters.sample_buff\[8\] _07554_ _07555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12833_ _04828_ _04838_ _04839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_69_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09818__A1 channels.freq2\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11625__A1 channels.pw2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_174_3604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12764_ _04765_ _04766_ _04769_ _04770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_56_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15552_ channels.sample2\[3\] _03220_ _07490_ _03344_ _07491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_174_3615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11715_ channels.sus_rel3\[2\] _03782_ _01278_ channels.sus_rel2\[2\] _03806_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_16_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14503_ _03374_ _06177_ _06500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15483_ _06891_ _06767_ _07427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12695_ _04478_ _04698_ _04700_ _04701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_56_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17222_ _00292_ clknet_leaf_93_clk channels.sample2\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_182_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11646_ _03737_ _03727_ _03739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_14434_ _06425_ _06430_ _06431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_108_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09046__A2 _01497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput14 bus_in[6] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17153_ _00223_ clknet_leaf_122_clk channels.freq3\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_142_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14365_ _05509_ _05774_ _06363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_181_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_103_clk clknet_5_13__leaf_clk clknet_leaf_103_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11577_ channels.freq3\[4\] _03688_ _03690_ _03691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_108_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08514__B _00129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16104_ _07978_ _07979_ _07980_ _07981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13316_ _05235_ _05238_ _05322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17084_ _00154_ clknet_leaf_108_clk channels.freq1\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10528_ _02733_ _02786_ _02787_ _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_123_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14296_ _06293_ _06294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_126_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16035_ _07880_ _07903_ _07914_ _07915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_13247_ _04470_ _04712_ _05253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10459_ _01164_ _02517_ _02720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_161_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13178_ _04742_ _05183_ _05184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__15347__B _06979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12129_ _04146_ _00514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_36_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16937_ _00016_ clknet_leaf_217_clk channels.lfsr\[3\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11166__I _03381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10070__I _02330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16868_ _00955_ _00956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_149_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15819_ _06897_ _07636_ _07711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_172_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16893__S _00975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16799_ _03490_ _01817_ _00882_ _00880_ _08462_ _08461_ _00904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai33_1
XFILLER_0_59_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09340_ _01013_ _01743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_177_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11616__A1 _03662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09080__B _01534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08475__I _01004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09271_ channels.lfsr\[2\]\[19\] _01701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11115__B _03333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14030__A2 _04341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_172_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12592__A2 _04597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14869__A1 filters.band\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_110_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08986_ _01435_ _01409_ _01448_ _01421_ _00065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10107__A1 _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15771__I _07663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08720__A1 _01201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09607_ _01875_ _01989_ _01990_ _01993_ _01994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_108_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09538_ _01927_ _01904_ _01905_ clk_trg\[1\] _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11607__A1 _03677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09276__A2 _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09469_ net2 _01787_ _01845_ _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__12280__A1 filters.res_lut\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15720__B _07333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11500_ _02324_ _03632_ _03636_ _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_152_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12480_ _04199_ _04485_ _04486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09028__A2 _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11431_ channels.accum\[1\]\[3\] _03593_ _03596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12635__I _04207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14150_ _06148_ _06017_ _06149_ _06150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_145_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11362_ _03554_ channels.adsr_state\[0\]\[1\] _03552_ _03555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__16849__A2 _03728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_130_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10594__A1 _02575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13101_ _05106_ _05107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10313_ _01156_ _02573_ _02574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14081_ _05987_ _05995_ _06081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_11293_ net8 _03499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__15521__A2 _07458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13032_ _05021_ _05028_ _05038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_10244_ _02504_ _02505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_167_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12370__I _04375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10175_ _02426_ _02405_ channels.pw3\[5\] _02436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__12099__A1 _01219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16777__I _02272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17771_ _00841_ clknet_leaf_205_clk channels.exp_periods\[2\]\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_128_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14983_ _06918_ _06954_ _00560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_128_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16722_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[7\] _08454_ _08451_ _08457_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13934_ _05803_ _05807_ _05936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_89_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16653_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[1\] _08267_ _08400_ _08401_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__15588__A2 _07518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13865_ _05865_ _05758_ _05866_ _05867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_159_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15604_ _01977_ _07538_ _07539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12816_ _03287_ _04197_ _04444_ _04822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_16584_ _08356_ _08360_ _00755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_158_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13796_ _05794_ _05798_ _05799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_57_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15535_ _03281_ _07463_ _07474_ _03375_ _07475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_173_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12747_ _04752_ _04753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_85_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15466_ _06875_ _07409_ _07411_ _07412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12678_ _04591_ _04678_ _04682_ _04683_ _04684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_84_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17205_ _00275_ clknet_leaf_174_clk channels.sample3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_11629_ channels.pw2\[6\] _03720_ _03722_ _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14417_ _06331_ _06345_ _06414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15397_ _07343_ _07348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17136_ _00206_ clknet_leaf_124_clk channels.atk_dec2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14348_ _06331_ _06345_ _06346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_25_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15856__I _01822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17067_ _00137_ clknet_leaf_104_clk filters.lp vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14279_ _06275_ _06277_ _06278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_100_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16018_ _07889_ _07895_ _07898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_90_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08840_ _01308_ _01311_ _01312_ _01159_ _01313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_97_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08771_ _01246_ _00052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_85_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11825__S _03886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_1_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16776__A1 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15579__A2 _03378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11624__I _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14251__A2 _06249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09323_ _01673_ _01734_ _01735_ _01677_ _00115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_177_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09254_ _01687_ _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_90_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_32_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09185_ channels.lfsr\[2\]\[6\] _01628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_32_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12565__A2 _04498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16700__A1 _08419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10328__A1 _02484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10879__A2 _02890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_145_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_145_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08969_ _01349_ _01432_ _01433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13817__A2 _05074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14865__I1 filters.band\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11828__A1 _01151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11980_ _03892_ _04053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_162_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10931_ channels.sample1\[2\] _03164_ _03166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_123_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13650_ _05527_ _05530_ _05654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10862_ _03031_ _02940_ _03114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_151_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_140_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12601_ _04604_ _04605_ _04607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_78_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13581_ _04176_ _05585_ _05586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10793_ _03019_ _03020_ _03046_ _03048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_66_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12532_ _04523_ _04524_ _04538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_15320_ _03468_ _06065_ _07278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_164_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12463_ _04279_ _04469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12365__I _04314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15251_ _01747_ channels.sample1\[11\] _07213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_151_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14202_ _06199_ _06200_ _06201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11414_ channels.accum\[2\]\[20\] _03586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_15182_ _07093_ _07094_ _07144_ _07145_ _07146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__14950__B1 channels.sample2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12394_ _04184_ _04400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_62_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_169_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_169_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14133_ _06128_ _06132_ _06133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_50_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11345_ _03096_ _03539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_105_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13505__A1 _05509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13505__B2 _05510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14064_ _06062_ _06064_ _06065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_11276_ _02334_ _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13015_ _05018_ _04515_ _05020_ _05021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_10227_ _01481_ _02487_ _02488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_123_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_182_3758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08932__A1 channels.freq3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_182_3769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10158_ _02406_ _02407_ _02419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_55_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17754_ _00824_ clknet_leaf_50_clk tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10089_ _02350_ _02351_ _02352_ _02354_ _00266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_14966_ _05647_ _06936_ _06937_ _06938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_16705_ tt_um_rejunity_sn76489.latch_control_reg\[0\] _08443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_13917_ _05834_ _05839_ _05919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_17685_ _00755_ clknet_5_11__leaf_clk tt_um_rejunity_sn76489.tone\[1\].gen.counter\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__16758__A1 _08453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14897_ filters.low\[28\] _06875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_18_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11444__I _01219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16636_ _01577_ _08388_ _08389_ _01702_ _00778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_13848_ _05850_ _05748_ _05851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_175_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16567_ _08344_ _08346_ _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_169_1304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13779_ _05769_ _05781_ _05782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_48_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15518_ filters.sample_buff\[0\] _07448_ _07451_ _07459_ _07460_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13992__A1 _04498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_23__f_clk_I clknet_3_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16498_ _08287_ _08288_ _00741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_128_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15449_ filters.low\[27\] _06862_ _07396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_26_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13744__A1 _05657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10558__A1 _02561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17119_ _00189_ clknet_leaf_115_clk channels.freq2\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_13_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09941_ channels.freq3\[9\] _02248_ _02243_ _02251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10523__I _01089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09872_ channels.ctrl_reg2\[4\] _02202_ _02199_ _02203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_230_clk_I clknet_5_17__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08823_ channels.ctrl_reg1\[1\] channels.sync_outs\[2\] _01295_ _01296_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_174_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08754_ _01232_ _01234_ _01235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09479__A2 _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_245_clk_I clknet_5_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12483__A1 _03413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08685_ channels.exp_counter\[0\]\[0\] channels.exp_counter\[1\]\[0\] channels.exp_counter\[2\]\[0\]
+ channels.exp_counter\[3\]\[0\] _01152_ _01168_ _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_174_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_68_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_156_Left_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_85_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09306_ _01721_ _01728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08663__I _01146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09651__A2 net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09237_ _01670_ _01671_ _01664_ _01672_ _01643_ _01644_ _01673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_8_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12185__I _04190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09168_ channels.lfsr\[3\]\[2\] _01614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14783__I0 filters.low\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09099_ _01300_ _01551_ _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XPHY_EDGE_ROW_165_Left_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11130_ _03191_ _03248_ _03197_ _03347_ _03348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XTAP_TAPCELL_ROW_147_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_147_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11061_ _03192_ _03283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_164_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10012_ channels.atk_dec3\[3\] _02292_ _02294_ _02300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12710__A2 _04714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14820_ _06795_ _06800_ _06805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_4_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15660__A1 channels.sample1\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14751_ _06741_ _06703_ _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11963_ _03903_ _03854_ _04032_ _04039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_59_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_174_Left_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11264__I _03473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13702_ _05612_ _05613_ _05706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_86_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10914_ _03154_ _03080_ _03155_ _00290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_17470_ _00540_ clknet_leaf_15_clk filters.band\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_168_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14682_ _04453_ _05883_ _06677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11894_ channels.env_vol\[0\]\[6\] _03965_ _03979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16421_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[12\] _08220_ _08227_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15412__B2 _07321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13633_ _05604_ _05637_ _05638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10845_ _03095_ _03097_ _03098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16352_ _08176_ _08177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08573__I _01089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13564_ _04630_ _05561_ _05569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10776_ _02955_ _03031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15303_ _03455_ _07244_ _07261_ _07262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_12515_ _04223_ _04232_ _04521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_16283_ net19 _07719_ _08140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13495_ _05500_ _05501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13726__A1 _03333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12446_ _04451_ _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15234_ _07176_ _07191_ _07196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_151_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12377_ _04334_ _04337_ _04382_ _04383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_15165_ _01761_ channels.sample2\[8\] _07130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11328_ _02103_ _03525_ _00334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14116_ _04740_ _04781_ _06116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15096_ _07035_ _07061_ _07063_ _00564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_120_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11439__I _02364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14151__A1 _05069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14047_ _05928_ _06046_ _06047_ _06048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_11259_ _03468_ _03226_ _03469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08905__A1 _01367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_173_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15998_ _07756_ _07751_ _07878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_167_Right_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_167_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17737_ _00807_ clknet_leaf_53_clk tt_um_rejunity_sn76489.control_tone_freq\[0\]\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14949_ _01759_ _01745_ channels.sample1\[0\] channels.sample2\[0\] _06922_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
Xclkbuf_leaf_74_clk clknet_5_9__leaf_clk clknet_leaf_74_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09330__A1 _01577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08470_ _00997_ net3 _00999_ _01000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_17668_ _00738_ clknet_leaf_80_clk tt_um_rejunity_sn76489.tone\[2\].gen.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_175_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_148_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16619_ _01638_ _08381_ _08383_ _01640_ _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_9_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12217__A1 _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_174_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17599_ _00669_ clknet_leaf_57_clk spi_dac_i.spi_dat_buff_0\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08483__I _01004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11440__A2 _03593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15706__A2 _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09022_ _01481_ _01482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_31_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_170_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09397__A1 _01742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09924_ _02154_ _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__15890__A1 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[2\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09855_ channels.pw2\[11\] _02191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10703__A1 _02710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_142_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08806_ _01278_ _01279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08658__I _01141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09786_ _02123_ _01898_ _02141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_1_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_134_Right_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12456__A1 _04448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08737_ channels.exp_counter\[1\]\[0\] _01105_ _01218_ _01220_ _01221_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11259__A2 _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_64_clk_I clknet_5_11__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08668_ _01151_ _01152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_120_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08599_ _01110_ _00016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_138_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10630_ _02886_ _02887_ _02888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_79_clk_I clknet_5_12__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09085__B1 _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_157_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10561_ _01689_ _02771_ _02821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11033__B _03256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_122_clk_I clknet_5_30__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11431__A2 _03593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12300_ _04285_ _04305_ _04306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_63_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13280_ _05267_ _05285_ _05286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_133_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_118_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10492_ _02750_ _02752_ _02753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_118_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12231_ _04236_ _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_32_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11814__S0 _03832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12162_ _04167_ _04168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_leaf_137_clk_I clknet_5_31__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11113_ _03331_ _03332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_9_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12093_ _04072_ _04104_ _04127_ _00497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16970_ _00049_ clknet_leaf_193_clk channels.exp_counter\[2\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15921_ _07800_ _07802_ _07795_ _07803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11044_ _03257_ _03258_ _03263_ _03267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_60_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09560__A1 channels.atk_dec1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15852_ _03735_ _07736_ _07737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_118_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15633__A1 channels.sample2\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14803_ _06769_ _06778_ _06789_ _06790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_15783_ _06791_ _07677_ _07686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_101_Right_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_56_clk clknet_5_8__leaf_clk clknet_leaf_56_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12995_ _04998_ _05000_ _05001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09312__A1 _01632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17522_ _00592_ clknet_leaf_21_clk filters.sample_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_169_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14734_ _06689_ _06726_ _06727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11946_ channels.env_counter\[2\]\[3\] _04013_ _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_169_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_177_3668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17453_ _00523_ clknet_leaf_191_clk channels.accum\[3\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12818__I _04780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14665_ _06537_ _06593_ _06660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11877_ _03539_ _03963_ _03964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11670__A2 _03759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16404_ _08213_ _08214_ _08211_ _00721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13947__A1 _04238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13616_ _03383_ _04342_ _04804_ _05621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_39_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17384_ _00454_ clknet_leaf_137_clk channels.env_counter\[2\]\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10828_ _03054_ _03080_ _03081_ _00278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14596_ _06563_ _06591_ _06592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_138_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16734__B _08459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16335_ channels.env_vol\[1\]\[5\] _08166_ _08168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13547_ _05439_ _05526_ _05552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10759_ _02882_ _03013_ _03014_ _00276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_41_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16266_ _07597_ _08129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13478_ _05308_ _05311_ _05483_ _05484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__09379__A1 _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13175__A2 _03470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15217_ _01772_ _02029_ _07160_ _07180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_129_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12429_ _04432_ _04426_ _04434_ _04435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_16197_ _08037_ _08051_ _08070_ _08071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_50_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12922__A2 _04927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15148_ _05416_ _07066_ _07114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_77_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10933__A1 channels.sample1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15079_ _07045_ _07046_ _07047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14675__A2 _05626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09551__A1 _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09640_ channels.sus_rel2\[5\] _01936_ _02001_ channels.freq2\[5\] _02026_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09571_ channels.freq1\[2\] _01954_ _01834_ channels.freq3\[10\] _01959_ _01960_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_78_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_47_clk clknet_5_10__leaf_clk clknet_leaf_47_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_117_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09303__A1 _01598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08522_ _01021_ _01035_ _01048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_65_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09005_ channels.freq3\[12\] _01079_ _01466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_143_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13166__A2 _05070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_76_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09907_ _02208_ _01869_ _02226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09838_ channels.freq2\[15\] _02171_ _02176_ _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11028__B _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09769_ channels.atk_dec1\[2\] _02126_ _02129_ _02130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_154_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_38_clk clknet_5_3__leaf_clk clknet_leaf_38_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11800_ _03890_ _03869_ _03838_ _03891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_139_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12780_ _04782_ _04785_ _04786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_159_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output27_I net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11731_ channels.atk_dec3\[7\] _01078_ _03780_ channels.atk_dec2\[7\] _03788_ channels.atk_dec1\[7\]
+ _03822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_51_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14450_ _06415_ _06446_ _06447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11662_ _03752_ _03753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13401_ _05406_ _04948_ _05407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10613_ _02768_ _02869_ _02871_ _02774_ _02872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_92_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11593_ channels.pw3\[2\] _03697_ _03698_ _03701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_36_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14381_ _06237_ _06377_ _06378_ _06379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_172_3576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16120_ _07960_ _07961_ _07959_ _07781_ _07997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__09947__I _02254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13332_ net69 _05336_ _05337_ _05338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10544_ _01687_ _02572_ _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16051_ _07853_ _07930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_133_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_133_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13263_ _04765_ _05268_ _05090_ _05269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10475_ _02566_ _02734_ _02735_ _02736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_51_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11168__A1 _03374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15002_ _03268_ _06947_ _06973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_150_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12214_ _04219_ _04220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13194_ _05154_ _05200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14106__A1 _06030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08584__A2 _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12145_ _04154_ _00522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_124_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15617__C _03395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12076_ channels.env_counter\[0\]\[7\] _04114_ _04118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16953_ _00032_ clknet_leaf_239_clk channels.lfsr\[3\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15904_ _07785_ _07786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11027_ filters.band\[1\] _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_95_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16884_ _01205_ _00955_ _00964_ _00968_ _00969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_21_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15606__A1 channels.sample2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_179_3708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15835_ _07721_ _07722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_29_clk clknet_5_0__leaf_clk clknet_leaf_29_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_91_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09631__B _01809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15766_ _03455_ _07670_ _07671_ _07674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12978_ _04972_ _04973_ _04984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_17505_ _00575_ clknet_leaf_249_clk filters.high\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14717_ _03422_ _06397_ _06711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11929_ _04011_ _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15697_ _07623_ _00605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17436_ _00506_ clknet_leaf_185_clk channels.accum\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14648_ _05509_ _06096_ _06643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_60_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15859__I _07741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14763__I _06752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17367_ _00437_ clknet_leaf_171_clk channels.pw2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14579_ _06420_ _06424_ _06575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_126_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16318_ _08156_ _00693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_166_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08761__I _01083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17298_ _00368_ clknet_leaf_186_clk channels.accum\[1\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_97_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14345__A1 _06337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16249_ filters.sample_buff\[4\] _08115_ _08117_ spi_dac_i.spi_dat_buff_0\[0\] spi_dac_i.spi_dat_buff_0\[1\]
+ _07728_ _08118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_42_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_58_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10906__A1 channels.sample2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09772__A1 channels.atk_dec1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10382__A2 _02555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12659__A1 _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09524__A1 channels.freq1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09524__B2 channels.ctrl_reg1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13320__A2 _04489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09623_ channels.ch3_env\[4\] _02009_ _01948_ channels.atk_dec1\[4\] _02010_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16270__A1 filters.sample_buff\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09554_ _01859_ _01943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09288__B1 _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13623__A3 _05624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08505_ _01008_ _01019_ _01032_ _01033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09485_ _01783_ _01836_ _01831_ _01876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__10437__A3 _02607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_154_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11398__A1 _03566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08671__I _01154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12193__I _04198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10260_ _01157_ _02520_ _02521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12898__A1 _04902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08566__A2 _01082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12921__I _04926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10191_ _02444_ _02445_ _02446_ _02452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__11570__A1 _03664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11537__I _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09515__A1 channels.sample3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09515__B2 clk_trg\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13950_ _04254_ _05185_ _05952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12901_ _04878_ _04891_ _04906_ _04907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_13881_ _05775_ _05883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_159_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15620_ _07552_ _07553_ _07554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_12832_ _04831_ _04833_ _04837_ _04838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_158_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15551_ _03297_ _07488_ _07489_ _03376_ _07490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_174_3605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12763_ _04709_ _04767_ _04768_ _04769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12822__A1 _04821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_174_3616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14502_ _06498_ _06499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_11714_ _03794_ _03805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_90_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15482_ _07416_ _07411_ _07425_ _07408_ _07418_ _07426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_12_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12694_ _04699_ _04697_ _04469_ _04696_ _04700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_83_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17221_ _00291_ clknet_leaf_94_clk channels.sample2\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_182_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14433_ _06428_ _06429_ _06430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_11645_ _03737_ _03728_ _03738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_52_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17152_ _00222_ clknet_leaf_143_clk channels.freq3\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput15 bus_in[7] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_14364_ _06359_ _05989_ _06362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12050__A2 _02354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11576_ _03689_ _03690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13199__I _05151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16103_ _07958_ _07968_ _07980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10061__A1 filters.cutoff_lut\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13315_ _05320_ _05305_ _05321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_17083_ _00153_ clknet_leaf_109_clk channels.freq1\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10527_ _02736_ _02782_ _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14295_ _06283_ _06293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_150_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16034_ _07908_ _07913_ _07914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_13246_ _05069_ _04750_ _05252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10458_ _02717_ _02718_ _02719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_58_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09754__A1 _01807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13177_ _04858_ _05183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10389_ _02627_ _02640_ _02649_ _02650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__10364__A2 _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15827__A1 _03194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12128_ channels.accum\[3\]\[12\] _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_36_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12059_ _04107_ _04108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09506__B2 channels.pw3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16936_ _00015_ clknet_leaf_216_clk channels.lfsr\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_53_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10116__A2 _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16867_ _00954_ _00955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14758__I _05546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15818_ _06882_ _07697_ _07709_ _07710_ _00639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_172_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16798_ _07759_ _00896_ _00903_ _00901_ _00819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_176_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15749_ _03374_ _07656_ _07657_ _07662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09270_ _01577_ _01589_ _01592_ _01700_ _00097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08493__A1 net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_99_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17419_ _00489_ clknet_leaf_139_clk channels.env_counter\[0\]\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09993__A1 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08796__A2 channels.ctrl_reg3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_9_clk clknet_5_5__leaf_clk clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_125_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_15__f_clk clknet_3_3_0_clk clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_141_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09745__A1 channels.ctrl_reg1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08985_ _01436_ _01446_ _01447_ _01448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_48_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11855__A2 _03934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16243__A1 _07924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09606_ channels.atk_dec3\[4\] _01991_ _01992_ channels.freq3\[12\] _01993_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__08666__I _01149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13057__A1 _04895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09537_ channels.sample3\[5\] _01927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_39_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09468_ _01000_ _01789_ _01859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08484__A1 filters.res_filt\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10291__A1 _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14557__A1 _05512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09399_ filters.mode_vol\[1\] _01794_ _01796_ _01797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11430_ _03595_ _03591_ _01348_ _03592_ _00366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_163_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09984__A1 _02252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11240__B1 _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11361_ _01585_ _03529_ _03531_ _03549_ _03554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_162_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_130_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10312_ channels.env_vol\[0\]\[6\] channels.env_vol\[1\]\[6\] _01142_ _02573_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13100_ filters.cutoff_lut\[16\] _04441_ _05106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11292_ _03497_ _03498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14080_ _05544_ _06080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_131_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10243_ _02503_ _02504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13031_ _04693_ _04992_ _05016_ _05036_ _05037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_167_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_167_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10174_ _01285_ _02435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_28_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11267__I _03476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17770_ _00840_ clknet_leaf_201_clk channels.exp_periods\[2\]\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14982_ filters.high\[2\] _06934_ _06951_ _06953_ _06954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_128_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16721_ _02298_ _08456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_13933_ _05918_ _05934_ _05935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_156_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16652_ _08399_ _08400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_159_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08576__I channels.clk_div\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13864_ _05750_ _05754_ _05866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_92_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_158_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15603_ _07513_ _07538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12815_ _04313_ _04820_ _04821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_9_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16583_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[6\] _08347_ _08358_ _08359_
+ _08360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_85_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13795_ _05795_ _05797_ _05798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_151_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15534_ channels.sample3\[2\] _07463_ _07474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12746_ _04751_ _04752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_139_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_127_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15465_ _07409_ _07410_ _07411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_13_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12677_ _04587_ _04590_ _04589_ _04683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_155_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17204_ _00274_ clknet_leaf_174_clk channels.sample3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14416_ _06316_ _06330_ _06413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11628_ _03673_ _03719_ _03724_ _00435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_142_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13071__I1 filters.band\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15396_ _07335_ _07347_ _06979_ _00580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_142_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10034__A1 _02314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17135_ _00205_ clknet_leaf_128_clk channels.atk_dec2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_163_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10346__I _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14347_ _06334_ _06344_ _06345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11559_ channels.freq2\[7\] _03670_ _03671_ _03678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_107_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17066_ _00136_ clknet_leaf_106_clk filters.mode_vol\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14278_ _06082_ _06163_ _06276_ _06277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_123_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16017_ _07896_ _07897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09727__A1 _02098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13229_ _04324_ _04405_ _05235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_90_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08770_ channels.exp_counter\[2\]\[3\] _01245_ _01235_ _01241_ _01246_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_16919_ _00966_ channels.exp_periods\[0\]\[2\] _00987_ _00990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_26_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_69_Left_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08486__I _01015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_177_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15821__B _07700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09322_ _01668_ _01734_ _01735_ _01671_ _00114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09663__B1 _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_168_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09253_ _01656_ _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12736__I _04198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11640__I _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_173_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09184_ _01621_ _01611_ _01625_ _01627_ _00084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_32_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13211__A1 _05211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_78_Left_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09966__A1 channels.pw3\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09281__I3 _01709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09718__A1 _01742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_149_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11525__A1 channels.pw1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10328__A2 _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08941__A2 _01360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08968_ _01430_ _01431_ _01432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09780__I _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_87_Left_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_162_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08899_ channels.accum\[0\]\[4\] channels.accum\[1\]\[4\] channels.accum\[2\]\[4\]
+ channels.accum\[3\]\[4\] _01146_ _01161_ _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XTAP_TAPCELL_ROW_162_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10930_ _03162_ _02831_ _03165_ _00296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_123_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15731__B _07648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10861_ _03088_ _02890_ _03113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_140_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12600_ _04604_ _04605_ _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_67_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13580_ _05504_ _05585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_109_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09654__B1 _01970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10792_ _03019_ _03020_ _03046_ _03047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_148_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10264__A1 _01482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12531_ filters.res_lut\[1\] _04168_ _04537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_82_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15250_ _01761_ channels.sample2\[11\] _07212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_164_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12462_ _04390_ _04468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_87_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09020__I _00010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15957__I _07722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14201_ _06115_ _06120_ _06200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09957__A1 _02240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11413_ _03578_ _01545_ _03585_ _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_152_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15181_ _07135_ _07138_ _07145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_12393_ _04200_ _04181_ _04399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_169_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14132_ _06129_ _06130_ _06131_ _06132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_169_3526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11344_ _03039_ _03536_ _03537_ _03538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_160_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09709__A1 channels.freq1\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13505__A2 _04758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14063_ _05877_ _05967_ net46 _06064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11275_ _03483_ _03484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11516__A1 _03513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_148_Right_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13014_ _04502_ _05019_ _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_123_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10226_ _02464_ _02466_ _02487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16788__I _00895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_182_3759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_242_clk clknet_5_18__leaf_clk clknet_leaf_242_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10157_ _02403_ _02417_ _02418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_17753_ _00823_ clknet_leaf_50_clk tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10088_ _02353_ _02354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_14965_ _01773_ channels.sample3\[0\] _06924_ _06937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_16704_ tt_um_rejunity_sn76489.latch_control_reg\[1\] _08442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_13916_ _05908_ _05917_ _05918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_17684_ _00754_ clknet_leaf_64_clk tt_um_rejunity_sn76489.tone\[1\].gen.counter\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14896_ _06856_ _06871_ _06872_ _06835_ _06873_ _06874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XTAP_TAPCELL_ROW_18_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16635_ _01698_ _08388_ _08389_ _01573_ _00777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_76_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15641__B _07573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13847_ _05743_ _05746_ _05850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16566_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[3\] _08345_ _08339_ _08346_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_57_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13778_ _05772_ _05780_ _05781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_48_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15517_ filters.sample_buff\[0\] _07458_ _07459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_57_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12556__I _04561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12729_ _04258_ _04485_ _04735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16497_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[3\] _08282_ _08252_ _08288_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13992__A2 _05990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15448_ filters.low\[27\] _07395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_26_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16930__A2 _00923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10007__A1 _02250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14771__I _06760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15379_ _03733_ _07332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_142_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17118_ _00188_ clknet_leaf_114_clk channels.freq2\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16899__S _00975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16694__A1 _08238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09940_ _02184_ _02250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_141_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17049_ _00119_ clknet_leaf_230_clk channels.lfsr\[1\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12291__I _04281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_115_Right_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09871_ _02193_ _02202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16446__A1 _04101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_233_clk clknet_5_17__leaf_clk clknet_leaf_233_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__15249__A2 channels.sample3\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08822_ _01294_ _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08753_ _01216_ _01233_ _01234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_75_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08684_ _01167_ _01168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_178_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13680__A1 _04512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12483__A2 _04488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_105_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13850__I _03376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08944__I _01257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09305_ _01615_ _01723_ _01727_ _01618_ _00105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10246__A1 _02484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12786__A3 _04444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09236_ channels.lfsr\[3\]\[12\] _01672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_174_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09939__A1 _02245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14932__A1 _06761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09167_ channels.lfsr\[1\]\[2\] _01613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_32_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09098_ _01548_ _01550_ _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__16685__A1 _08419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_147_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11060_ filters.low\[3\] _03282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10011_ _02298_ _02299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_224_clk clknet_5_20__leaf_clk clknet_leaf_224_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08914__A2 _01360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_125_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14750_ _06739_ _03222_ _06740_ _06741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_169_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11962_ _04027_ _04037_ _04038_ _00455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13701_ _05616_ _05636_ _05704_ _05705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_86_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10913_ channels.sample2\[7\] _03150_ _03155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14681_ _06332_ _05980_ _06571_ _06676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11682__B1 _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11893_ _03128_ _03977_ _03978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_98_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16420_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[11\] _08223_ _08226_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13632_ _05616_ _05636_ _05637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10844_ _03096_ _02940_ _03071_ _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_6_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16351_ _02356_ _03937_ _08176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11434__B1 _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13563_ _05566_ _05567_ _05568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_6_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10775_ _02624_ _02994_ _03030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15302_ _05968_ _07245_ _07261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12514_ _04431_ _04519_ _04520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16282_ _08138_ _08139_ _07740_ _00674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_125_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13494_ _05351_ _05500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_180_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15233_ _03410_ _07064_ _07195_ _07089_ _00569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_152_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12445_ _04450_ _04451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_22_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15164_ _01770_ channels.sample3\[8\] _07129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_151_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12376_ _04335_ _04336_ _04382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14115_ _06109_ _06114_ _06115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_11327_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[0\] _03522_ _03524_ _03525_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15095_ filters.high\[6\] _07062_ _06775_ _07063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14046_ _04752_ _05828_ _05721_ _05930_ _06047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__14151__A2 _05350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11258_ filters.low\[15\] _03468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_215_clk clknet_5_21__leaf_clk clknet_leaf_215_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10209_ channels.pw2\[3\] _02470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08905__A2 _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11189_ filters.sample_filtered\[10\] _03403_ _03404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_15997_ _07748_ _07874_ _07876_ _07877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_17736_ _00806_ clknet_leaf_63_clk tt_um_rejunity_sn76489.control_tone_freq\[0\]\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14948_ _04431_ _04519_ _06920_ _06921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_0_82_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10476__A1 _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17667_ _00737_ clknet_leaf_47_clk net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14879_ _06851_ _06858_ _06859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__16600__A1 tt_um_rejunity_sn76489.chan\[1\].attenuation.in vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16618_ _01632_ _08381_ _08383_ _01635_ _00766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_17598_ _00668_ clknet_leaf_58_clk spi_dac_i.spi_dat_buff_0\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16549_ _08326_ _08330_ _08331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_175_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12286__I _04291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08841__A1 _01304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09021_ channels.accum\[0\]\[13\] channels.accum\[1\]\[13\] channels.accum\[2\]\[13\]
+ channels.accum\[3\]\[13\] _01138_ _01480_ _01481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_116_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14914__A1 _06889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_143_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10951__A2 _03136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09923_ _02234_ _02235_ _02237_ _00217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12153__A1 _04158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_206_clk clknet_5_22__leaf_clk clknet_leaf_206_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09854_ _02188_ _02181_ _02190_ _00195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08805_ _01277_ _01278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_142_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09785_ _01819_ _02133_ _02140_ _00176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15642__A2 _07568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08736_ _01219_ _01220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08667_ _01150_ _01151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13580__I _05504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_71_Right_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_166_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08598_ channels.lfsr\[3\]\[3\] _01110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_165_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10219__A1 _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_154_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_157_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10560_ _01550_ _02567_ _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_64_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11033__C _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13708__A2 _04924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09219_ _01652_ _01634_ _01657_ _01651_ _00089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10491_ _01158_ _02581_ _02751_ _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_118_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12230_ _04235_ _04236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_121_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11814__S1 _01171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12392__A1 _04265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_80_Right_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_121_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12161_ _04166_ _04167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_31_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_15_Left_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10942__A2 _03052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11112_ _03247_ _03248_ _03250_ _03330_ _03331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XTAP_TAPCELL_ROW_9_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12092_ channels.env_counter\[0\]\[14\] _04107_ _04127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15456__B _07333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15920_ _07784_ _07797_ _07801_ _07798_ _07802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_11043_ _03242_ _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08849__I _01320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15851_ _07721_ _07733_ _07734_ _07730_ _07735_ _07736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_14802_ _06780_ _06781_ _06779_ _06789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_118_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15782_ _07681_ _07685_ _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12994_ _04969_ _04999_ _04965_ _05000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__13644__A1 _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17521_ _00591_ clknet_leaf_18_clk filters.sample_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14733_ _03440_ _03222_ _06725_ _06726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_11945_ _04009_ _04023_ _04024_ _04025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_93_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17452_ _00522_ clknet_leaf_157_clk channels.accum\[3\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14664_ _06594_ _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_177_3669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11876_ _03961_ _03947_ _03962_ _03963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16403_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[7\] _08209_ _08214_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13615_ _03364_ _04854_ _05220_ _05620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__11407__B1 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17383_ _00453_ clknet_leaf_136_clk channels.env_counter\[2\]\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_145_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13947__A2 _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10827_ _01977_ _02975_ _03081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14595_ _06590_ _06591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_54_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16334_ _03964_ _08165_ _08167_ _00698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15149__A1 _03345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13546_ _05439_ _05526_ _05551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08823__A1 channels.ctrl_reg1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10758_ _01927_ _02975_ _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16972__CLK clknet_5_23__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17549__D _00619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16265_ _08121_ _08128_ _00668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13477_ _05309_ _05310_ _05483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_82_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10689_ _02908_ _02911_ _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_15216_ _07152_ _07177_ _07178_ _07179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12428_ _04419_ _04433_ _04434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_113_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16196_ _08049_ _08050_ _08070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_129_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_244_clk_I clknet_5_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15147_ _07098_ _07112_ _07113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_168_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12359_ _04319_ _04327_ _04365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_168_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15321__A1 filters.low\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15078_ _01745_ channels.sample1\[5\] _07046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14029_ _06028_ _05925_ _06029_ _06030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__13883__A1 _05440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10697__A1 _02555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09570_ _01955_ _01957_ _01958_ _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_175_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08521_ _01027_ _01036_ _01029_ _01047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17719_ _00789_ clknet_leaf_62_clk tt_um_rejunity_sn76489.tone\[0\].gen.counter\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_65_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09067__A1 _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12744__I _04489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09004_ _01464_ _01465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10924__A2 _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13575__I _05514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09906_ _02160_ _02219_ _02225_ _00212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_6_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08669__I _00010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09837_ _02157_ _02170_ _02177_ _00191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__16812__B2 _01817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09768_ _02093_ _02129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13626__A1 _03316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08719_ _01179_ channels.exp_periods\[3\]\[3\] _01203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_179_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09699_ _01767_ _02074_ _02079_ _00151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11823__I _03905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_159_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11730_ _01292_ _03820_ _03791_ _03821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_84_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11044__B _03263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11661_ _03096_ _03540_ _03752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_154_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13400_ _04940_ _05406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_92_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10612_ _02402_ _02770_ _02870_ _02871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_135_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14380_ _06238_ _06239_ _06378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_137_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11592_ _03662_ _03696_ _03700_ _00423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_172_3577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13331_ _05234_ _05239_ _05337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10612__A1 _02402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10543_ _02712_ _02802_ _02803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_52_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16050_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[2\] _07927_ _07928_
+ _07760_ _07878_ _07929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_126_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13262_ _05092_ _05268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_133_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_23_Left_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10474_ _02611_ _02651_ _02735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15001_ _06939_ _05035_ _06972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11168__A2 _03378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12213_ _04218_ _04219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__13686__S _05179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13193_ _05138_ _05152_ _05199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12144_ channels.accum\[3\]\[20\] _04154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_103_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12075_ _04037_ _04113_ _04117_ _00489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16952_ _00031_ clknet_leaf_239_clk channels.lfsr\[3\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15903_ _07784_ tt_um_rejunity_sn76489.chan\[0\].attenuation.in _07785_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11026_ _03249_ _03250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_95_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16883_ _00944_ _00960_ _00968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__16803__A1 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[0\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15606__A2 _03395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15834_ _07717_ _07721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_179_3709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_32_Left_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12977_ _04981_ _04982_ _04983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15765_ _06737_ _07664_ _07673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17504_ _00574_ clknet_leaf_248_clk filters.high\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11928_ _01581_ _04005_ _01102_ _04011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_14716_ _06067_ _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15696_ channels.exp_periods\[3\]\[0\] _07623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09203__I _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14647_ _06553_ _06554_ _06641_ _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_17435_ _00505_ clknet_leaf_178_clk channels.accum\[3\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09049__A1 _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11859_ channels.env_vol\[0\]\[1\] _03942_ _03949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_60_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17366_ _00436_ clknet_leaf_101_clk channels.pw2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14578_ _06565_ _06573_ _06574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_166_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16317_ channels.env_counter\[3\]\[14\] _08156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_126_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13529_ _05534_ _03346_ _05535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17297_ _00367_ clknet_leaf_178_clk channels.accum\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_41_Left_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_141_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16248_ _08116_ _08117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_63_clk_I clknet_5_11__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10084__I clk_trg\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16179_ spi_dac_i.spi_dat_buff_1\[6\] _07729_ _07869_ spi_dac_i.spi_dat_buff_1\[7\]
+ _03734_ _08054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_58_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_78_clk_I clknet_5_12__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_50_Left_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_177_1267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_121_clk_I clknet_5_27__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09622_ _01877_ _02009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_37_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09553_ channels.pw1\[10\] _01890_ _01941_ channels.ctrl_reg1\[2\] _01942_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09288__B2 _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08504_ _01010_ _01032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__13623__A4 _05626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09484_ _01874_ _01875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12292__B1 _04296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_136_clk_I clknet_5_31__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_114_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14033__A1 _04750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_154_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_154_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12898__A2 _04903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10190_ _02447_ _02450_ _02451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_30_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15836__A2 _04776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13847__A1 _05743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09515__A2 _01904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09071__S0 _01139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12900_ _04895_ _04900_ _04905_ _04906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_13880_ _05782_ _05880_ _05881_ _05882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_119_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12831_ _04834_ _04835_ _04836_ _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__13075__A2 _04758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15550_ channels.sample3\[3\] _07453_ _07489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_167_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12762_ _04714_ _04715_ _04768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_51_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_174_3606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12822__A2 _04827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_174_3617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14501_ _06494_ _06497_ _06498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11713_ _03794_ _03803_ _03804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_56_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15481_ _07412_ _07419_ _07425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_56_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12693_ _04255_ _04699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_37_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09958__I _02254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14432_ _04802_ _05448_ _06429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17220_ _00290_ clknet_leaf_173_clk channels.sample2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11644_ _01264_ _03737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_108_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17151_ _00221_ clknet_leaf_143_clk channels.freq3\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_142_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14363_ _06243_ _06244_ _06360_ _06361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xinput16 bus_we net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_135_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11575_ _02333_ _03689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08885__S0 _01308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16102_ _07958_ _07968_ _07979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13314_ _05313_ _05319_ _05320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_91_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_181_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17082_ _00152_ clknet_leaf_106_clk channels.freq1\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10526_ _02736_ _02782_ _02786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14294_ _03347_ _06080_ _06292_ _06187_ _00533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_123_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12338__A1 _03316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16033_ _07820_ _07904_ _07912_ _07913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13245_ _04228_ _04740_ _05251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10457_ _02681_ _02682_ _02702_ _02718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_161_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13176_ _05181_ _04537_ _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_62_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_107_Left_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10388_ _02643_ _02648_ _02649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_62_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11561__A2 _01871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12127_ _04145_ _00513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12058_ _04106_ _04107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16935_ _00014_ clknet_leaf_216_clk channels.lfsr\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_53_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11009_ _03233_ _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_5_17__f_clk_I clknet_3_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16866_ _03544_ _03755_ _00953_ _00952_ _00954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_15817_ _02353_ _07710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_172_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16797_ net11 _00897_ _00903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14263__A1 _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11463__I _01104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17516__CLK clknet_5_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15748_ _06506_ _07652_ _07661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_142_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14015__A1 _04259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09690__A1 _01781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15679_ filters.sample_buff\[13\] _07448_ _07608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_99_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17418_ _00488_ clknet_leaf_138_clk channels.env_counter\[0\]\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_16_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17349_ _00419_ clknet_leaf_100_clk channels.freq3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15515__A1 channels.sample1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_110_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11638__I _03731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15818__A2 _07697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08984_ _01438_ _01431_ _01445_ _01447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_177_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09108__I _01460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16491__A2 _08282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12501__A1 _04504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12501__B2 _04506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09605_ _01833_ _01992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09536_ channels.sus_rel1\[1\] _01899_ _01901_ channels.atk_dec1\[1\] _01926_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11068__A1 filters.high\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09467_ channels.freq1\[0\] _01855_ _01857_ channels.ctrl_reg1\[0\] _01858_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_176_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08484__A2 _01013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14006__A1 _04742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08682__I _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14557__A2 _05796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15754__A1 _03394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09398_ _01752_ _01796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_129_Right_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_73_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11240__A1 _03243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11360_ _03553_ _00338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_132_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_130_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10311_ _02519_ channels.env_vol\[3\]\[6\] _02571_ _02572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_85_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11291_ _03490_ _03491_ _03492_ _03496_ _03497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_85_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13030_ _05035_ _05031_ _05036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_10242_ channels.env_vol\[0\]\[0\] channels.env_vol\[1\]\[0\] channels.ch3_env\[0\]
+ channels.env_vol\[3\]\[0\] _01145_ _01159_ _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_30_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_167_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10173_ channels.pw1\[5\] _02434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_167_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14981_ _06935_ _06950_ _06952_ _06953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13763__I _05671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16720_ _08453_ _08446_ _08455_ _00796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13932_ _05920_ _05933_ _05934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_57_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16651_ _08398_ _08399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13863_ _05750_ _05755_ _05865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_18_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14245__A1 _04697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15602_ filters.sample_buff\[6\] _07529_ _07537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_12814_ _04819_ _04820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16582_ _08353_ _08357_ _08301_ _08359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13794_ _04487_ _05796_ _05797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15533_ _07462_ _07469_ _07473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12745_ _04750_ _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_5_21__f_clk clknet_3_5_0_clk clknet_5_21__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_57_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15464_ filters.low\[28\] _06717_ _07410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_72_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12676_ _04677_ _04674_ _04675_ _04681_ _04682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_167_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12559__A1 _03317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14415_ _06410_ _06411_ _06412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17203_ _00273_ clknet_leaf_179_clk channels.sample3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_182_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11627_ channels.pw2\[5\] _03720_ _03722_ _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_170_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15395_ _07062_ _07346_ _07347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_154_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17134_ _00204_ clknet_leaf_127_clk channels.ctrl_reg2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_14346_ _06343_ _06344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09975__A2 _01881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11558_ _01817_ _03677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17065_ _00135_ clknet_leaf_106_clk filters.mode_vol\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10509_ _02541_ _02770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_14277_ _06085_ _06162_ _06276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11489_ _03511_ _03625_ _03629_ _00391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_122_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16016_ _07889_ _07895_ _07896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_100_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13228_ _05148_ _05232_ _05233_ _05234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_55_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10362__I _02622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13159_ _05138_ _05152_ _05164_ _05165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_176_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11298__A1 _02314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16918_ _00989_ _00853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16849_ _01581_ _03728_ _01087_ _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__14787__A2 _04160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09321_ _01730_ _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09663__A1 filters.res_filt\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09663__B2 channels.sample3\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09252_ channels.lfsr\[3\]\[14\] _01686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_91_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09183_ _01626_ _01627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13211__A2 _05216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_181_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09966__A2 _02266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12970__A1 _04448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12752__I _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_rebuffer11_I _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11368__I _02974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08967_ _01423_ _01419_ _01429_ _01431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__11289__A1 net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08677__I _01160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08898_ _01365_ _01366_ _01367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_162_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_123_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10860_ _03087_ _03110_ _03111_ _03112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_123_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09519_ _01873_ _01889_ _01907_ net22 _01909_ _01910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_91_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09654__A1 channels.sus_rel3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10791_ _03044_ _03045_ _03046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09654__B2 channels.freq1\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12530_ _04535_ _04171_ _04536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_136_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11461__A1 _03612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12461_ _04254_ _04467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_151_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14200_ _06109_ _06198_ _06199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11412_ channels.accum\[2\]\[19\] _03556_ _03585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11213__A1 _03422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15180_ _07113_ _07117_ _07144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_12392_ _04265_ _04397_ _04398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14950__A2 channels.sample1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14131_ _04367_ _05347_ _06131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_169_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11343_ _02707_ _02711_ _03537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_104_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14062_ _05966_ _05963_ _06063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_11274_ _02088_ _01849_ _03483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_39_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13013_ _04497_ _04515_ _05019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10225_ _02476_ _02477_ _02451_ _02485_ _02486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_33_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10156_ _02414_ _02416_ _02417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_146_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13269__A2 _05268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14466__A1 _05510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17752_ _00822_ clknet_leaf_48_clk tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10087_ _01724_ _02353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14964_ _06922_ _06923_ _06925_ _06936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16703_ tt_um_rejunity_sn76489.latch_control_reg\[2\] _08441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_57_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13915_ _05912_ _05916_ _05917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_17683_ _00753_ clknet_leaf_66_clk tt_um_rejunity_sn76489.tone\[1\].gen.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14895_ _06853_ _06863_ _06718_ _06873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_89_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16634_ _01694_ _08388_ _08389_ _01695_ _00776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_57_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13846_ _05846_ _05848_ _05849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_134_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16565_ _08243_ _08345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09645__A1 channels.ch3_env\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13777_ _05773_ _05779_ _05780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10989_ _03204_ _03214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_174_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09645__B2 channels.atk_dec1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11452__A1 _03600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15516_ _07456_ _07457_ _07458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_128_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12728_ _04253_ _04179_ _04734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16496_ _08285_ _08286_ _08287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_128_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09211__I _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15447_ _07382_ _07394_ _00584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12659_ _04322_ _04633_ _04634_ _04615_ _04665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__15194__A2 channels.sample2\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15378_ _07326_ _07329_ _07330_ _07331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_108_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12952__A1 _04701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17117_ _00187_ clknet_leaf_115_clk channels.freq2\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__12572__I _04525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14329_ _04806_ _05280_ _06327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17048_ _00118_ clknet_5_17__leaf_clk channels.lfsr\[1\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15883__I tt_um_rejunity_sn76489.chan\[1\].attenuation.in vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10092__I _01082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09870_ _02193_ _02201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_96_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09881__I _01779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08821_ _01293_ _01294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09008__S0 _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08752_ _01186_ _01231_ _01199_ _01233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08497__I _01015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16928__B _02272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08683_ _01166_ _01167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_174_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13680__A2 _04447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15551__C _03376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11651__I _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09304_ _01608_ _01723_ _01727_ _01613_ _00104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10246__A2 _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09235_ channels.lfsr\[1\]\[12\] _01671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_57_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10267__I _02527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13196__A1 _05138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09166_ channels.lfsr\[0\]\[2\] _01612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09097_ _01549_ _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_160_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14696__A1 _03412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_164_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10010_ _01775_ _02298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__16437__A2 _08238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09999_ _02289_ _01867_ _02290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_125_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14999__A2 _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13120__A1 _05122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09324__B1 _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11961_ channels.env_counter\[2\]\[6\] _04030_ _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09875__A1 _02155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13700_ _05618_ _05635_ _05704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10912_ _02365_ _03154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14680_ filters.band\[30\] _04633_ _06675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11682__B2 _03766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11892_ _03976_ _03542_ _03946_ _03977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13631_ _05618_ _05635_ _05636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10843_ _02961_ _03096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_168_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12226__A3 _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14620__A1 _06614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13562_ _05497_ _05523_ _05567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16350_ _08175_ _00706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10774_ _03028_ _02840_ _03029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11434__B2 _03592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_181_Right_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12513_ _04435_ _04518_ _04519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_15301_ filters.low\[15\] _06065_ _07260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_16281_ spi_dac_i.spi_dat_buff_1\[11\] _08117_ _08139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14872__I _06706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13493_ _05323_ net47 _05498_ _05499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_137_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_180_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12444_ _04375_ _04450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_43_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15232_ _07192_ _07193_ _07194_ _07195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_63_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12934__A1 _04844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15163_ _07127_ _07128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12375_ _04365_ _04380_ _04381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__10905__I _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14114_ _06112_ _06113_ _06114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_105_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11326_ _01740_ _03523_ _03524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15094_ _06982_ _07062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_14045_ _04929_ _05465_ _05930_ _05828_ _06046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_11257_ filters.high\[15\] _03467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_120_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10208_ _02463_ _02467_ _02468_ _02469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11188_ _03399_ _03402_ _03403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10139_ channels.pw1\[10\] _01285_ _02400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15996_ _07841_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[0\] _07746_
+ _07876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_17735_ _00805_ clknet_leaf_63_clk tt_um_rejunity_sn76489.control_tone_freq\[1\]\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14947_ _04558_ _04690_ _04691_ _06920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_106_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17666_ _00736_ clknet_leaf_41_clk tt_um_rejunity_sn76489.noise\[0\].gen.counter\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14878_ _06854_ _06857_ _06858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_16617_ _01625_ _08381_ _08383_ _01629_ _00765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_15_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09618__A1 channels.pw1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13829_ _05829_ _05830_ _05831_ _05832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_174_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17597_ _00667_ clknet_leaf_40_clk spi_dac_i.spi_dat_buff_0\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12217__A3 _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14611__A1 _06298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09618__B2 channels.ctrl_reg1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16548_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[1\] _08267_ _08329_ _08330_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_35_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11425__B2 _03592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10087__I _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16479_ _08266_ _08271_ _08272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_143_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_151_clk clknet_5_29__leaf_clk clknet_leaf_151_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_5_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13178__A1 _04742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09020_ _00010_ _01480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_182_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08780__I _01253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09922_ channels.sus_rel2\[4\] _02236_ _02232_ _02237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12153__A2 _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09853_ channels.pw2\[10\] _02182_ _02189_ _02190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_142_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08804_ _01276_ _01277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09784_ channels.atk_dec1\[7\] _02134_ _02138_ _02140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13102__A1 _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08735_ _01100_ _01219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_1_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08666_ _01149_ _01150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_139_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08597_ _01109_ _00015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_157_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_142_clk clknet_5_30__leaf_clk clknet_leaf_142_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__16355__A1 channels.ch3_env\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13169__A1 _05069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09218_ _01653_ _01654_ _01646_ _01655_ _01142_ _01656_ _01657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_106_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10490_ _01688_ _02580_ _02751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_118_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11719__A2 _03809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12916__A1 _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09149_ channels.lfsr\[3\]\[0\] _01597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_135_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13101__I _05106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12392__A2 _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12160_ _03189_ _03181_ _03195_ _04166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__10242__I2 channels.ch3_env\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11111_ filters.band\[6\] _03330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_12091_ _04068_ _04104_ _04126_ _00496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_9_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11042_ _03244_ _03265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10155__A1 _01566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15850_ spi_dac_i.counter\[2\] _07735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14801_ _06706_ _06787_ _06788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__09848__A1 channels.pw2\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15781_ filters.low\[18\] _07682_ _07684_ _07685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12993_ _04211_ _04966_ _04999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13644__A2 _03376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17520_ _00590_ clknet_leaf_18_clk filters.sample_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14732_ _03439_ _06710_ _06725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11944_ _03833_ _04015_ _03888_ _04024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_87_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17451_ _00521_ clknet_leaf_158_clk channels.accum\[3\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11875_ _03538_ _03951_ _03962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14663_ _06656_ _06657_ _06658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16402_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[6\] _08212_ _08213_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13614_ _04864_ _04445_ _05619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10826_ _03057_ _03079_ _03080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_67_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17382_ _00452_ clknet_leaf_129_clk channels.env_counter\[2\]\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14594_ _06574_ _06589_ _06590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_55_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16333_ channels.env_vol\[1\]\[4\] _08166_ _08167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_171_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10757_ _02979_ _03012_ _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_13545_ net35 net39 _05531_ _05550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_133_clk clknet_5_31__leaf_clk clknet_leaf_133_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09481__C1 _01871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_164_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16264_ filters.sample_buff\[9\] _08125_ _08122_ spi_dac_i.spi_dat_buff_0\[5\] spi_dac_i.spi_dat_buff_0\[6\]
+ _08127_ _08128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_13476_ _05478_ _05481_ _05482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_152_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10688_ _02909_ _02910_ _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_153_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12907__A1 _04833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12427_ _04415_ _04426_ _04433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_15215_ _07156_ _07161_ _07178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_16195_ _08058_ _08059_ _08068_ _08069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_124_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08587__A1 _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12358_ _04328_ _04363_ _04364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_51_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15146_ filters.low\[8\] _07111_ _07112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_11_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11309_ _03506_ _03508_ _03510_ _02273_ _00330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_15077_ _01759_ channels.sample2\[5\] _07045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12289_ _04294_ _04295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_120_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14028_ _04290_ _04397_ _05732_ _06027_ _06029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__09000__A2 _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10697__A2 _02638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14777__I _06765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09839__A1 _02160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15979_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[1\] _07856_ _07859_
+ _07771_ _07860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_179_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_175_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08520_ _01046_ _00001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_17718_ _00788_ clknet_leaf_62_clk tt_um_rejunity_sn76489.tone\[0\].gen.counter\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_17649_ _00719_ clknet_leaf_50_clk tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_82_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_124_clk clknet_5_27__leaf_clk clknet_leaf_124_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_144_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09003_ _01453_ _01454_ _01464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08578__A1 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13571__A1 _05568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_83_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12760__I _04753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09905_ channels.atk_dec2\[7\] _02220_ _02224_ _02225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09836_ channels.freq2\[14\] _02171_ _02176_ _02177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11309__C _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09767_ _02110_ _02125_ _02128_ _00170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_154_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13626__A2 _04163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17572__CLK clknet_5_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08718_ channels.exp_periods\[2\]\[3\] _01202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09698_ channels.freq1\[10\] _02075_ _02077_ _02079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_2__f_clk clknet_3_0_0_clk clknet_5_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_159_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08649_ _01135_ _00041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_139_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11660_ _03746_ _03750_ _03751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_83_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09058__A2 _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10611_ _01705_ _02771_ _02870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_154_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_115_clk clknet_5_26__leaf_clk clknet_leaf_115_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11591_ channels.pw3\[1\] _03697_ _03698_ _03700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_172_3567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13330_ _05234_ _05239_ _05336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_88_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_172_3578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10542_ _01157_ _02635_ _02801_ _02802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_135_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13261_ _05198_ _05266_ _05267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10473_ _02611_ _02651_ _02734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_33_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12212_ filters.cutoff_lut\[6\] filters.res_lut\[6\] _04217_ _04218_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15000_ net37 _06969_ _06970_ _06971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_62_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13192_ _05166_ _05191_ _05197_ _05198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12143_ _04153_ _00521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13314__A1 _05313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12074_ channels.env_counter\[0\]\[6\] _04114_ _04117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16951_ _00030_ clknet_leaf_224_clk channels.lfsr\[3\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15902_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[2\] _07784_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_11025_ filters.filter_step\[0\] _03249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_16882_ _00967_ _00839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15833_ spi_dac_i.counter\[0\] _07720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13617__A2 _05621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11628__A1 _03673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15764_ _07669_ _07672_ _00623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12976_ _04811_ _04812_ _04982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14290__A2 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17503_ _00573_ clknet_leaf_21_clk filters.high\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14715_ _06298_ _06698_ _06705_ _06708_ _06709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_11927_ _03880_ _04009_ _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_169_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15695_ _07615_ _07484_ _07622_ _07269_ _00604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__10300__A1 _01328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17434_ _00504_ clknet_leaf_187_clk channels.accum\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14646_ _04576_ _06383_ _06555_ _06641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11858_ _03944_ _03947_ _03948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09049__A2 _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_106_clk clknet_5_15__leaf_clk clknet_leaf_106_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__12053__A1 _04101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10809_ _03029_ _03035_ _03033_ _03063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16319__A1 _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17365_ _00435_ clknet_5_25__leaf_clk channels.pw2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11789_ _03879_ _03880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14577_ _06567_ _06572_ _06573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_144_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16316_ _08155_ _00692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_172_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13528_ filters.low\[0\] _05534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_153_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17296_ _00366_ clknet_leaf_186_clk channels.accum\[1\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_141_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16247_ _07720_ _07717_ _08116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_97_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13459_ _05229_ _05465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_97_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16178_ _08033_ _08036_ _08052_ _08053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_141_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15377__B _07240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_58_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15129_ _07093_ _07094_ _07095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_75_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10119__A1 channels.ctrl_reg1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09621_ filters.res_filt\[4\] _02007_ _01939_ channels.sample3\[8\] _02008_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__11924__I _04006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13608__A2 _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09552_ _01857_ _01941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11619__A1 channels.pw2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08503_ _01009_ _00129_ _01031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09483_ net7 _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11145__B _03361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12292__B2 _04297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_93_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14033__A2 _04884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15781__A2 _07682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13792__A1 _04200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10275__I _02535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13544__A1 _05527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10358__A1 _01534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08971__A1 _01422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15836__A3 _07722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13847__A2 _05746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09071__S1 _01480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09819_ _02105_ _02163_ _02165_ _00185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09732__C _02103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16797__A1 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12830_ _04473_ _04377_ _04836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_243_clk_I clknet_5_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12761_ _04714_ _04715_ _04767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_68_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_174_3607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14500_ _06304_ _06395_ _06496_ _06497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_174_3618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11712_ _03802_ _03803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15480_ filters.high\[30\] _06919_ _07424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12692_ _04694_ _04281_ _04696_ _04697_ _04698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__15221__A1 _01762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11643_ _03728_ _03736_ _00438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14431_ _06426_ _06427_ _06428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_154_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17150_ _00220_ clknet_leaf_142_clk channels.sus_rel2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_11574_ _03679_ _03688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14362_ _06359_ _05891_ _06245_ _06360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xinput17 rst net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__10141__S0 _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16101_ _07956_ _07978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08885__S1 _01160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13313_ _05317_ _05318_ _05319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10525_ _02359_ _02783_ _02785_ _00271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_17081_ _00151_ clknet_leaf_107_clk channels.freq1\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14293_ _05975_ _06291_ _06292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_24_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16032_ _07910_ _07911_ _07912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13244_ _05174_ _05248_ _05249_ _05250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_165_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10456_ _02709_ _02715_ _02716_ _02717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_122_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13175_ filters.high\[16\] _03470_ _05180_ _05181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_27_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10387_ _02646_ _02647_ _02648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_20_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08962__A1 channels.freq2\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12126_ channels.accum\[3\]\[11\] _04145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08962__B2 channels.freq1\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12057_ _01319_ _04004_ _01032_ _04106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_16934_ _00013_ clknet_leaf_215_clk channels.lfsr\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_53_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11008_ _03232_ _03233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16865_ _01267_ _02455_ channels.clk_div\[0\] _01094_ _00953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_15816_ _06888_ _07698_ _07709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16796_ _07755_ _00896_ _00902_ _00901_ _00818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_88_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14263__A2 _06261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15747_ _07659_ _07660_ _00618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_133_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12959_ _04512_ _04420_ _04965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15678_ _07598_ _07607_ _00602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_23_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15212__A1 _03394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09690__A2 _01970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17417_ _00487_ clknet_leaf_135_clk channels.env_counter\[0\]\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14629_ _06578_ _06579_ _06624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_16_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15763__A2 _07670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17348_ _00418_ clknet_leaf_101_clk channels.freq3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16491__B _08252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17279_ _00349_ clknet_leaf_163_clk channels.accum\[2\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09884__I _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_1308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_73_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08983_ _01438_ _01431_ _01445_ _01446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_11_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16779__A1 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10512__A1 _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11654__I _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09604_ _01866_ _01991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_155_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_108_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16666__B _08292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_108_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09535_ filters.mode_vol\[1\] _01791_ _01896_ channels.pw3\[1\] _01925_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_39_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09130__A1 _01577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09466_ _01856_ _01789_ _01853_ _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_65_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14006__A2 _05588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15203__A1 _03374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09397_ _01742_ _01793_ _01795_ _00133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_136_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13765__A1 _05563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10579__A1 _02687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10310_ _02518_ _02570_ _02571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11290_ _03495_ _03496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_105_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10241_ _02501_ _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_113_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10172_ _02425_ _02429_ _02431_ _02433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_TAPCELL_ROW_167_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_167_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_121_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14980_ _06907_ _06952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_13931_ _05927_ _05932_ _05933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_16650_ _08393_ _08398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_5_9__f_clk_I clknet_3_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_182_clk_I clknet_5_19__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13862_ _05852_ _05855_ _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_9_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16576__B _08301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15601_ filters.sample_buff\[7\] _07484_ _07536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12813_ _04818_ _04819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12256__A1 filters.res_lut\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16581_ _08353_ _08357_ _08358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_clkbuf_leaf_62_clk_I clknet_5_11__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13793_ filters.high\[23\] filters.band\[23\] _03187_ _05796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09121__A1 _01300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15532_ filters.sample_buff\[1\] _07468_ _07472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12744_ _04489_ _04750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_96_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_197_clk_I clknet_5_23__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15463_ _07395_ _06766_ _07409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__12395__I _04400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12675_ _04592_ _04679_ _04680_ _04681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_182_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17202_ _00272_ clknet_leaf_179_clk channels.sample3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14414_ _06347_ _06370_ _06411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12559__A2 _04506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13756__A1 _05547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11626_ _03668_ _03719_ _03723_ _00434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_25_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_77_clk_I clknet_5_12__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15394_ _07342_ _07345_ _07346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_108_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17133_ _00203_ clknet_leaf_117_clk channels.ctrl_reg2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_170_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14345_ _06337_ _06342_ _06343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11557_ _03675_ _03669_ _03676_ _00412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_94_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_94_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17064_ _00134_ clknet_leaf_105_clk filters.mode_vol\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10508_ _01542_ _02539_ _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11488_ channels.freq1\[1\] _03626_ _03627_ _03629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_123_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14276_ _06189_ _06192_ _06274_ _06275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_0_100_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16015_ _07773_ _07891_ _07894_ _07895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_123_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10439_ _02677_ _02678_ _02700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13227_ _04280_ _05231_ _04825_ _05230_ _05233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_55_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_135_clk_I clknet_5_31__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13158_ _05154_ _05157_ _05163_ _05164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_20_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17573__D _00643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12109_ _04136_ _00504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13089_ _05094_ _05095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_85_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_15_clk_I clknet_5_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16917_ _00962_ channels.exp_periods\[0\]\[1\] _00987_ _00989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16848_ _08419_ _00936_ _00836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_137_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16779_ net10 _00886_ _00890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09320_ _01728_ _01734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09251_ channels.lfsr\[1\]\[14\] _01685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_103_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09182_ _01588_ _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_149_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08958__I _01321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08966_ _01423_ _01419_ _01429_ _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__11289__A2 _03494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12486__A1 _04487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08897_ channels.freq2\[4\] _01275_ _01288_ channels.freq1\[4\] _01366_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__09351__A1 _01748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_95_clk clknet_5_13__leaf_clk clknet_leaf_95_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_162_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_162_Right_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_168_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12238__A1 _03273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_123_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09518_ _01908_ _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_149_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12789__A2 _04314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10790_ _03021_ _03022_ _03043_ _03045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_TAPCELL_ROW_140_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09654__A2 _01943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11333__B _03517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09449_ _00997_ _01784_ _00999_ _01840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_137_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12460_ _04319_ _04327_ _04380_ _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_75_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11411_ _03584_ _03581_ _01539_ _03582_ _00358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_12391_ _04396_ _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_117_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14130_ _04371_ _05185_ _06130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11342_ _02710_ _03536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_169_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_169_3528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11273_ _03243_ _03481_ _03482_ _03245_ _03466_ _00322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_14061_ _06059_ _06061_ _06062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__08917__A1 _01377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13012_ _04497_ _05018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10224_ _02432_ _02480_ _02485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09590__A1 channels.ctrl_reg1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09590__B2 _01977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10155_ _01566_ _02415_ _02409_ _02404_ _02416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_100_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17751_ _00821_ clknet_leaf_48_clk tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10086_ net8 _02351_ _02352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14963_ _06928_ _06930_ _06935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_leaf_86_clk clknet_5_12__leaf_clk clknet_leaf_86_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_16702_ _07798_ _08437_ _08440_ _00793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13914_ _05913_ _05914_ _05915_ _05916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_17682_ _00752_ clknet_leaf_70_clk tt_um_rejunity_sn76489.tone\[1\].gen.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14894_ _06855_ _06871_ _06872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_16633_ _08382_ _08389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_18_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13845_ _05660_ _05742_ _05847_ _05848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_18_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16564_ _08342_ _08343_ _08344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_58_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13776_ _05777_ _05778_ _05779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_97_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10988_ _03208_ _03211_ _03179_ _03213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_168_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15515_ channels.sample1\[0\] _03400_ _07457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12727_ _04228_ _04272_ _04733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16495_ _08277_ _08284_ _08244_ _08286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_167_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13729__A1 _03350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15446_ filters.high\[26\] _06934_ _07391_ _07393_ _07394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12658_ _04639_ _04640_ _04646_ _04650_ _04664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_170_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11609_ _01780_ _01848_ _03711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__12401__A1 _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15377_ _07326_ _07329_ _07240_ _07330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12589_ _04594_ _04171_ _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_17116_ _00186_ clknet_leaf_111_clk channels.freq2\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14328_ _05909_ _05092_ _06326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17047_ _00117_ clknet_leaf_238_clk channels.lfsr\[1\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14259_ _06142_ _06157_ _06258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08908__B2 channels.freq1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08820_ _01292_ _01293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09581__A1 channels.ch3_env\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09581__B2 channels.pw1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09008__S1 _01154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14457__A2 _05446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08751_ _01186_ _01199_ _01231_ _01232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_174_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_77_clk clknet_5_12__leaf_clk clknet_leaf_77_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_40_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09333__A1 _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08682_ _01165_ _01166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_139_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_105_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_68_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13968__A1 _05969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09636__A2 _02019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09303_ _01598_ _01723_ _01727_ _01602_ _00103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_152_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09234_ channels.lfsr\[0\]\[12\] _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_125_Left_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09165_ _01610_ _01611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14393__A1 _06192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09096_ channels.accum\[0\]\[20\] channels.accum\[1\]\[20\] channels.accum\[2\]\[20\]
+ channels.accum\[3\]\[20\] _01138_ _01153_ _01549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_142_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14145__A1 filters.band\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14696__A2 _03378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10706__A1 _02676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_134_Left_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08688__I _01171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09998_ _01779_ _02289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15645__A1 channels.sample2\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_181_3750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08949_ _01412_ _01413_ _01414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_125_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_68_clk clknet_5_11__leaf_clk clknet_leaf_68_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_4_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11960_ _04019_ _04036_ _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_4_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10911_ _03147_ _03052_ _03153_ _00289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11682__A2 _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11891_ _03961_ _03753_ _03976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13630_ _05623_ _05634_ _05635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10842_ _03063_ _03070_ _03095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11063__B _03284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13561_ _05499_ _05522_ _05566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12631__A1 _03256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_143_Left_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_137_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10773_ _02602_ _03028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_149_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15300_ _06918_ _07259_ _00572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12512_ _04438_ _04517_ _04518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_16280_ net20 _07719_ _08138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13492_ _05324_ _05222_ _05329_ _05498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_124_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15231_ _07192_ _07193_ _07086_ _07194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_164_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12443_ _04372_ _04449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_63_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_43_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15162_ _07107_ _07108_ _07126_ _07127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12374_ _04370_ _04373_ _04379_ _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_105_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10193__I channels.pw2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14136__A1 _06105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14113_ _04711_ _04817_ _06113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11325_ _03521_ _03523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_50_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15093_ _07037_ _07060_ _07061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_127_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11256_ filters.sample_filtered\[15\] _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14044_ _05913_ _06043_ _06044_ _06045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_152_Left_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10207_ _02464_ _02466_ _01481_ _02468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_24_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11187_ filters.high\[10\] _03401_ _03402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11370__A1 _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10138_ _02389_ _02390_ channels.pw3\[10\] _02399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_89_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15995_ _07874_ _07875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xclkbuf_leaf_59_clk clknet_5_8__leaf_clk clknet_leaf_59_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_17734_ _00804_ clknet_leaf_63_clk tt_um_rejunity_sn76489.control_tone_freq\[1\]\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10069_ _02330_ _02340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14946_ _06908_ _06919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_82_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17665_ _00735_ clknet_leaf_57_clk tt_um_rejunity_sn76489.noise\[0\].gen.counter\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12848__I _04271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14877_ net32 _06855_ _06856_ _06857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__10476__A3 _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16616_ _01620_ _08381_ _08383_ _01622_ _00764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_13828_ _04753_ _05466_ _05831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_161_Left_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_17596_ _00666_ clknet_leaf_39_clk spi_dac_i.spi_dat_buff_0\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__16764__B _00877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16547_ _08328_ _08329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13759_ _05666_ _05677_ _05761_ _05762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_63_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16478_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[1\] _08267_ _08270_ _08271_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_127_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15429_ _07373_ _07374_ _07377_ _07378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12925__A2 _04928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10936__A1 channels.sample1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_170_Left_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09892__I _02174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09921_ _02226_ _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_106_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_146_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09852_ _02175_ _02189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11361__A1 _01585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08803_ _01275_ _01276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11148__B _03364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09783_ _01814_ _02133_ _02139_ _00175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_142_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13102__A2 _04215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08734_ _01169_ _01217_ _01218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_1_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08665_ _01148_ _01149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12861__A1 _04852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12758__I _04211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08596_ channels.lfsr\[3\]\[2\] _01109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09132__I _01082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_157_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09217_ _01155_ _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14366__A1 _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09148_ channels.lfsr\[1\]\[0\] _01596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_162_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_135_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09079_ _01533_ _01534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11110_ filters.low\[6\] _03329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_12090_ channels.env_counter\[0\]\[13\] _04107_ _04126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_9_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11041_ filters.sample_filtered\[2\] _03264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11352__A1 _03534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09307__I _01728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15618__A1 channels.sample2\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14800_ filters.low\[19\] filters.band\[19\] _06755_ _06787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_157_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09751__B _02113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15780_ _07683_ _07684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_118_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12992_ _04465_ _04495_ _04997_ _04998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_118_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14841__A2 _03473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14731_ net30 _06721_ _06723_ _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11943_ _03833_ _03888_ _04015_ _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_54_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16043__A1 _07838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17450_ _00520_ clknet_leaf_195_clk channels.accum\[3\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14662_ _06523_ _06533_ _06657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11874_ _03751_ _03961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_86_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16594__A2 _08274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16401_ _08191_ _08212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_54_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13613_ _05482_ _05490_ _05617_ _05618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_32_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17381_ _00451_ clknet_leaf_134_clk channels.env_counter\[2\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_157_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10825_ _03078_ _03079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14883__I _06706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14593_ _06576_ _06580_ _06588_ _06589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_27_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16332_ _08159_ _08166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_67_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13544_ _05527_ _05530_ _05549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_109_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_125_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10756_ _02982_ _03011_ _03012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_82_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09481__C2 channels.freq3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08823__A3 _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13499__I _05504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16263_ _07727_ _08127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13475_ _05479_ _05480_ _05481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_54_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10687_ _02914_ _02925_ _02943_ _02944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_54_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15214_ _07156_ _07161_ _07177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_140_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12907__A2 _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12426_ _04415_ _04432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_113_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16194_ _08064_ _08067_ _08068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_153_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10918__A1 channels.sample2\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14832__B _06765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09784__A1 channels.atk_dec1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08587__A2 _01100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15145_ _07101_ _07105_ _07110_ _07111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_105_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11040__B1 _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16603__I _08374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12357_ _04348_ _04351_ _04363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_168_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11591__A1 channels.pw3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11308_ _03499_ _03509_ _03510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15076_ _01769_ channels.sample3\[5\] _07044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12288_ _04198_ _04294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11718__I0 channels.atk_dec1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09536__B2 channels.atk_dec1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14027_ _04397_ _05732_ _06027_ _04290_ _06028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_11239_ _03450_ _03451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10146__A2 channels.pw2\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11343__A1 _02707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09217__I _01155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15978_ _07780_ _07858_ _07859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13096__A1 _04886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_165_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17717_ _00787_ clknet_leaf_67_clk tt_um_rejunity_sn76489.tone\[0\].gen.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14929_ filters.low\[31\] filters.band\[31\] _03477_ _06904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_26_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12843__A1 _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12843__B2 _04848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17648_ _00718_ clknet_leaf_50_clk tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_82_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17579_ _00649_ clknet_leaf_34_clk spi_dac_i.counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09472__B1 _01862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14899__A2 _03476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09002_ channels.accum\[0\]\[12\] _01463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_115_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13020__A1 _04996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08578__A2 _01093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11582__A1 _03675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_113_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09527__A1 _01762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11657__I _02687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09904_ _02216_ _02224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_6_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09527__B2 channels.pw2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11334__A1 _03515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09835_ _02175_ _02176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09766_ channels.atk_dec1\[1\] _02126_ _02120_ _02128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13087__A1 _04764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13626__A3 _05208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08717_ _01176_ _01201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_69_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09697_ _01757_ _02074_ _02078_ _00150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xrebuffer40 _05228_ net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_69_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08648_ channels.env_vol\[3\]\[5\] _01135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_96_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15799__I _07663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08579_ _01092_ _01094_ _01095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_25_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10610_ _01556_ _02567_ _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11590_ _03639_ _03696_ _03699_ _00422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_137_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_137_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10073__A1 _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_172_3568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10541_ _02529_ _02634_ _02801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_172_3579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13260_ _05203_ _05241_ _05265_ _05266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_10472_ _02652_ _02673_ _02732_ _02733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_161_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09766__A1 channels.atk_dec1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12211_ _04166_ _04217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_103_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13191_ _05134_ _05165_ _05197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12142_ channels.accum\[3\]\[19\] _04153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14511__A1 _03380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12073_ _04034_ _04113_ _04116_ _00488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16950_ _00029_ clknet_leaf_239_clk channels.lfsr\[3\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15901_ _07767_ _07771_ _07782_ _07783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11024_ _03193_ _03248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_16881_ _00966_ channels.exp_periods\[2\]\[2\] _00937_ _00967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_21_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15832_ _07718_ _07719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15763_ _03439_ _07670_ _07671_ _07672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12975_ _04978_ _04979_ _04980_ _04981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_59_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14714_ _06693_ _06707_ _06702_ _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_99_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17502_ _00572_ clknet_leaf_14_clk filters.high\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11926_ _03935_ _04009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15694_ _07619_ _07621_ _07622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14027__B1 _06027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09129__S0 _01201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17433_ _00503_ clknet_leaf_182_clk channels.accum\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_170_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14645_ _06472_ _04576_ _06640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_170_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11857_ _03946_ _03947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_60_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10808_ _02961_ _02939_ _03062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17364_ _00434_ clknet_leaf_171_clk channels.pw2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_14576_ _06568_ _06571_ _06572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_83_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11788_ channels.env_counter\[0\]\[0\] channels.env_counter\[1\]\[0\] channels.env_counter\[2\]\[0\]
+ channels.env_counter\[3\]\[0\] _01151_ _01167_ _03879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_172_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16315_ channels.env_counter\[3\]\[13\] _08155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10064__A1 _02314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13527_ _05532_ _05533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_166_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10739_ _02502_ _02994_ _02995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17295_ _00365_ clknet_leaf_182_clk channels.accum\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16246_ _07741_ _08115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13458_ _05326_ _05462_ _05463_ _05464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_24_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09757__A1 _01814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12409_ _04414_ _04351_ _04415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_16177_ _08037_ _08051_ _08052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_23_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13389_ _05129_ _05130_ _05395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_88_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_58_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15128_ _07026_ _07036_ _07060_ _07082_ _07094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_142_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15059_ _07026_ _07027_ _07028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10119__A2 _01286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09620_ _01844_ _02007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_71_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09551_ _01773_ _01002_ _01790_ filters.mode_vol\[2\] _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08502_ _01026_ _01030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09482_ _01835_ _01843_ _01865_ _01872_ _01873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_53_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15230__A2 _07168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_175_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10055__A1 _02289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09996__A1 channels.ctrl_reg3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09748__A1 _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13544__A2 _05530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_132_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15049__A2 channels.sample3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09818_ channels.freq2\[8\] _02164_ _02158_ _02165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09749_ _02106_ _02116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12760_ _04753_ _04766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_9_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13480__A1 _04278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output25_I net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_174_3608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11711_ _03801_ _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_174_3619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12691_ _04392_ _04697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_90_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15221__A2 channels.sample2\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14430_ _04805_ _05187_ _06427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11642_ channels.clk_div\[0\] _03732_ _03735_ _03736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_154_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09320__I _01728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14361_ _04575_ _06359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11573_ _03679_ _03687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16100_ _07954_ _07975_ _07976_ _07977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_24_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10141__S1 _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13312_ _05315_ _05316_ _05314_ _05318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_107_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17080_ _00150_ clknet_leaf_107_clk channels.freq1\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10524_ channels.sample3\[0\] _02784_ _02785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15478__B _07333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14292_ _06286_ _06290_ _06291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_108_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16031_ _07813_ _07822_ _07911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13243_ _04255_ _04392_ _04405_ _04751_ _05249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_21_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12338__A3 _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10455_ _02699_ _02700_ _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_33_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13174_ filters.band\[16\] _05179_ _05180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10386_ _02509_ _02594_ _02513_ _02647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_131_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12125_ _04144_ _00512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_92_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_176_Right_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12056_ _04104_ _04105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16933_ _00012_ clknet_leaf_193_clk channels.ring_outs\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_53_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09911__A1 _02179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11007_ _03231_ _03232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16864_ _00947_ _00949_ _00951_ _00952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_74_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15815_ _06875_ _07697_ _07708_ _07269_ _00638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_16795_ net10 _00897_ _00902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15746_ _03360_ _07656_ _07657_ _07660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08478__A1 filters.res_filt\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12958_ _04963_ _04964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13471__A1 _05313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11909_ _03991_ _03992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15677_ filters.sample_buff\[12\] _07447_ _07523_ _07606_ _07607_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_114_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12889_ _04834_ _04892_ _04894_ _04895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_158_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15212__A2 _07162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17416_ _00486_ clknet_leaf_131_clk channels.env_counter\[0\]\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14628_ _05909_ _05561_ _06623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_16_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10037__A1 _02316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17347_ _00417_ clknet_leaf_100_clk channels.freq3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14559_ _06553_ _06554_ _06555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_126_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_5_26__f_clk_I clknet_3_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17278_ _00348_ clknet_leaf_153_clk channels.accum\[2\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_141_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16229_ _08077_ _08092_ _08100_ _08101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12591__I _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08982_ _01444_ _01445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_143_Right_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09902__A1 channels.atk_dec2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09405__I _01017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09603_ channels.sus_rel3\[4\] _01963_ _01887_ channels.freq1\[12\] _01990_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_79_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_108_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09534_ channels.pw1\[9\] _01891_ _01893_ channels.freq2\[9\] _01924_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08469__A1 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09666__B1 _01899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09465_ _00997_ net3 _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__11473__B1 _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15203__A2 _07133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09396_ filters.mode_vol\[0\] _01794_ _01763_ _01795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09140__I _01588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09969__A1 _02252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10579__A2 _02777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11528__A1 _02326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10240_ _02500_ _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_132_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10171_ _01541_ _02425_ _02429_ _02431_ _02432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_112_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_167_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_167_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_110_Right_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13930_ _05928_ _05929_ _05931_ _05932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__09315__I _01730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13861_ _03284_ _05545_ _05863_ _05653_ _00529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_69_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15600_ _07498_ _07535_ _00596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12812_ _04817_ _04818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_69_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16580_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[6\] _08328_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[6\]
+ _08357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13792_ _04200_ _05500_ _05795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15531_ _07382_ _07471_ _00591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_57_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12743_ _04748_ _04749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_96_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15462_ _07389_ _07404_ _07405_ _07362_ _07407_ _07408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_182_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12674_ _04608_ _04609_ _04680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08880__A1 _01341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17201_ _00271_ clknet_leaf_169_clk channels.sample3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_155_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14413_ _06314_ _06346_ _06410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11625_ channels.pw2\[4\] _03720_ _03722_ _03723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14953__A1 _05647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15393_ _07343_ _07344_ _07345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_108_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17132_ _00202_ clknet_leaf_117_clk channels.ctrl_reg2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09275__I3 _01704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14344_ _06338_ _06341_ _06342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_11556_ channels.freq2\[6\] _03670_ _03671_ _03676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_94_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17063_ _00133_ clknet_leaf_105_clk filters.mode_vol\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10507_ _02538_ _02768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_94_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14275_ _06253_ _06273_ _06274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11487_ _02308_ _03625_ _03628_ _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_122_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16014_ _07773_ _07892_ _07893_ _07894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_123_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13226_ _04280_ _05229_ _05230_ _05231_ _05232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10438_ _02697_ _02698_ _02699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_0_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_55_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12192__A1 filters.res_lut\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_245_clk clknet_5_0__leaf_clk clknet_leaf_245_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13157_ _05159_ _05162_ _05163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XPHY_EDGE_ROW_29_Left_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10369_ _02543_ _02630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_104_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12108_ channels.accum\[3\]\[2\] _04136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13088_ _05087_ _05090_ _05093_ _05094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_174_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12039_ _04061_ _04090_ _04095_ _00475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16916_ _00988_ _00852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12495__A2 _04500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16847_ tt_um_rejunity_sn76489.clk_counter\[4\] _00935_ _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_178_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15433__A2 _06910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13444__A1 _05446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16778_ _07821_ _00885_ _00888_ _00889_ _00813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_87_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15729_ _07646_ _07647_ _00613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_87_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_38_Left_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09250_ channels.lfsr\[0\]\[14\] _01684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_103_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09181_ _01622_ _01623_ _01616_ _01624_ _01605_ _01607_ _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_172_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16697__A1 _08242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10981__A2 _03205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_47_Left_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_242_clk_I clknet_5_18__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_236_clk clknet_5_16__leaf_clk clknet_leaf_236_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_149_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_149_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08965_ _01427_ _01428_ _01429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_166_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08896_ channels.freq3\[4\] _01075_ _01365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_127_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13435__A1 _05440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10249__A1 _01497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09517_ _01874_ _01908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09448_ _01786_ net1 _01839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_13_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09379_ _01777_ _01743_ _01778_ _00128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_19_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11410_ channels.accum\[2\]\[18\] _03584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_46_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12390_ _04395_ _04396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_34_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11341_ _02805_ _03535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_127_1230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_169_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_3529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14060_ _05879_ _05962_ _06060_ _06061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_11272_ _03465_ _03480_ _03482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__15756__B _07648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_227_clk clknet_5_17__leaf_clk clknet_leaf_227_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13011_ _05011_ _05012_ _05004_ _05017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_63_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10223_ _02395_ _02418_ _02424_ _02483_ _02484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XANTENNA__11921__A1 _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09590__A2 _01941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10154_ _02398_ _02399_ _02400_ _02415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_100_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17750_ _00820_ clknet_leaf_47_clk tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14962_ _06908_ _06934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10085_ _02088_ _01905_ _02351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_55_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16701_ _07798_ _08437_ _08318_ _08440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13913_ _04317_ _04927_ _05915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17681_ _00751_ clknet_leaf_69_clk tt_um_rejunity_sn76489.tone\[1\].gen.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14893_ _06854_ _06864_ _06871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_89_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13790__I _05690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16632_ _08380_ _08388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13844_ _05662_ _05741_ _05847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_18_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13426__A1 _05423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16563_ _08336_ _08341_ _08292_ _08343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13775_ _04764_ _05775_ _05778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10987_ _03179_ _03208_ _03211_ _03212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_174_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_48_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_1308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12726_ _04706_ _04730_ _04731_ _04732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_48_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15514_ channels.sample2\[0\] _06066_ _07455_ _03344_ _07456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_16494_ _08277_ _08284_ _08285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08853__A1 channels.freq3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15445_ _06909_ _07392_ _07393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14926__A1 _06720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13729__A2 _04192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10660__A1 _02662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12657_ _04655_ _04657_ _04659_ _04663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_182_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11608_ _01740_ _03710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_25_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15376_ _07327_ _06754_ _07328_ _07329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__12401__A2 _04406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12588_ _04593_ _04594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_81_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17115_ _00185_ clknet_leaf_111_clk channels.freq2\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14327_ _06319_ _06324_ _06325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_53_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11539_ _03662_ _03658_ _03663_ _00407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17046_ _00116_ clknet_leaf_236_clk channels.lfsr\[1\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14258_ _06255_ _06256_ _06257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__14154__A2 _05588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15351__A1 _07295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15666__B _07573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12165__A1 filters.res_lut\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_218_clk clknet_5_21__leaf_clk clknet_leaf_218_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13209_ _05213_ _05214_ _05215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_111_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14189_ _06091_ _06099_ _06188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_110_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11912__A1 _01584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08750_ _01222_ _01231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_144_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12468__A2 _04471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16497__B _08252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08681_ _01164_ _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_136_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_85_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09302_ _01580_ _01723_ _01727_ _01596_ _00102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_158_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12640__A2 _04645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09233_ channels.lfsr\[2\]\[13\] _01669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_35_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10651__A1 _02657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_173_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15420__I filters.high\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09164_ _01590_ _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_161_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10564__I _02823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09095_ _01537_ _01543_ _01548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_181_clk_I clknet_5_19__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14145__A2 _04186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_209_clk clknet_5_17__leaf_clk clknet_leaf_209_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__15893__A2 tt_um_rejunity_sn76489.chan\[1\].attenuation.in vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_61_clk_I clknet_5_9__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11903__A1 _03905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_164_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12171__A4 filters.high\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09997_ _02242_ _02282_ _02288_ _00240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_196_clk_I clknet_5_23__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_181_3740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_3751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08948_ channels.freq2\[8\] _01277_ _01289_ channels.freq1\[8\] _01413_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_125_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_76_clk_I clknet_5_14__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09324__A2 _01734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08879_ _01299_ _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_99_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10910_ channels.sample2\[6\] _03150_ _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11890_ _03960_ _03974_ _03975_ _00446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_169_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10841_ _03091_ _03093_ _03094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_94_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13560_ _05562_ _05564_ _05565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_149_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10772_ _02995_ _02996_ _03026_ _03027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_66_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12631__A2 _04566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_134_clk_I clknet_5_31__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12511_ _04440_ _04496_ _04516_ _04517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_164_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13491_ _05346_ _05354_ _05496_ _05497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_82_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15230_ _07164_ _07168_ _07170_ _07193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_14_clk_I clknet_5_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12442_ _04353_ _04447_ _04448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_35_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_43_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15161_ _01771_ _01977_ _07109_ _07126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_105_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12373_ _04312_ _04378_ _04379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_149_clk_I clknet_5_31__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14112_ _06110_ _06111_ _06112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_11324_ _03521_ _03522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14136__A2 _06135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15092_ _07055_ _07059_ _07060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_105_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_29_clk_I clknet_5_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14043_ _05914_ _05915_ _06044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11255_ _03452_ _03460_ _03464_ _03465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_120_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10206_ _01481_ _02464_ _02466_ _02467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11186_ _03400_ _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15636__A2 _07568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10137_ _02397_ _01250_ channels.pw2\[10\] _02398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13647__A1 _05547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15994_ _07750_ _07754_ _07874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_17733_ _00803_ clknet_leaf_64_clk tt_um_rejunity_sn76489.control_tone_freq\[1\]\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10068_ _02299_ _02331_ _02339_ _00260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14945_ _01932_ _06918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15505__I _07446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17664_ _00734_ clknet_leaf_57_clk tt_um_rejunity_sn76489.noise\[0\].gen.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14876_ _06839_ _06846_ _06718_ _06856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_134_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16615_ _08382_ _08383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10881__A1 _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13827_ _04864_ _05721_ _05830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17595_ _00665_ clknet_leaf_39_clk spi_dac_i.spi_dat_buff_0\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_147_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16546_ _08327_ _08328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13758_ _05669_ _05676_ _05761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_58_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16349__B1 _01334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12709_ _04274_ _04295_ _04715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10633__A1 _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16477_ _08269_ _08270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13689_ _05688_ _05692_ _05693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_171_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15572__A1 filters.sample_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15428_ _07374_ _07376_ _07377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_182_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11189__A2 _03403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10384__I _02590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15359_ filters.low\[19\] _06499_ _07313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08685__S0 _01152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15396__B _06979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09920_ _02226_ _02235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09003__A1 _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17029_ _00006_ clknet_leaf_240_clk filters.res_lut\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_180_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08789__I _01261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_146_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09851_ _02187_ _02188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__16824__A1 _01776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08802_ _01274_ _01275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11361__A2 _03529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09782_ channels.atk_dec1\[6\] _02134_ _02138_ _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13638__A1 _05553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08733_ _01216_ _01217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08664_ _01147_ _01148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_68_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09413__I _01806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_120_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08595_ _01108_ _00014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14063__A1 _05877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16246__I _07741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_157_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_91_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09216_ channels.lfsr\[3\]\[9\] _01655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16690__B _01753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09147_ channels.lfsr\[0\]\[0\] _01595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_162_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_118_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10927__A2 _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_135_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09078_ channels.accum\[0\]\[18\] channels.accum\[1\]\[18\] channels.accum\[2\]\[18\]
+ channels.accum\[3\]\[18\] _01495_ _01496_ _01533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_124_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11040_ _03243_ _03261_ _03262_ _03245_ _03263_ _00308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__11352__A2 _03544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13629__A1 _05629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12991_ _04466_ _04494_ _04997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_118_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11942_ _04008_ _04021_ _04022_ _00451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14730_ _06722_ _06712_ _06723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16865__B channels.clk_div\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14661_ _06526_ _06532_ _06656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11873_ _03938_ _03960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16400_ _08208_ _08210_ _08211_ _00720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_129_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13612_ _05484_ _05489_ _05617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10824_ _03047_ _03077_ _03078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_17380_ _00450_ clknet_leaf_132_clk channels.env_counter\[2\]\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14592_ _06583_ _06587_ _06588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_45_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13801__A1 _04705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16331_ _08157_ _08165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13543_ _05533_ _05535_ _05536_ _05548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_94_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10755_ _02983_ _03010_ _03011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_39_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_153_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09481__B2 channels.sus_rel2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10091__A2 _02351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16262_ _08121_ _08126_ _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13474_ _03364_ _04854_ _04804_ _05480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_36_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10686_ _02896_ _02913_ _02943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_70_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15213_ _05533_ _07174_ _07175_ _07176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_12425_ _04309_ _04429_ _04430_ _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_16193_ _08065_ _08066_ _08067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_129_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10918__A2 _03156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15144_ _07106_ _07109_ _07110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11040__A1 _03243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12356_ _04310_ _04360_ _04361_ _04362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__11040__B2 _03263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11307_ _03507_ _03509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15075_ _07018_ _07041_ _07042_ _07043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12287_ _04187_ _04293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_121_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11718__I1 channels.sus_rel1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14026_ _05625_ _06027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09536__A2 _01899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11238_ filters.sample_filtered\[13\] _03450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11343__A2 _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15609__A2 _07543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_27__f_clk clknet_3_6_0_clk clknet_5_27__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11169_ _03373_ _03231_ _03384_ _03385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_101_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15977_ _07772_ _07857_ _07858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13096__A2 _04890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17716_ _00786_ clknet_leaf_73_clk tt_um_rejunity_sn76489.tone\[0\].gen.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_171_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14928_ _06901_ _06896_ _06902_ _06903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_136_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12843__A2 _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17647_ _00717_ clknet_leaf_50_clk tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14045__A1 _04929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14859_ _06835_ _06840_ _06841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_82_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17578_ _00648_ clknet_leaf_34_clk spi_dac_i.counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_11_Left_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16529_ _08135_ _08314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_156_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12594__I _04296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09472__A1 channels.sus_rel3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09472__B2 channels.pw2\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09001_ _01422_ _01459_ _01462_ _00066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12359__A1 _04319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10909__A2 _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11938__I _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09903_ _02157_ _02219_ _02223_ _00211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09527__A2 _01844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_130_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10137__A3 channels.pw2\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12531__A1 filters.res_lut\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09834_ _02174_ _02175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09765_ _02105_ _02125_ _02127_ _00169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13087__A2 _05092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08716_ channels.exp_periods\[0\]\[3\] channels.exp_periods\[1\]\[3\] _01187_ _01200_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11098__A1 _03310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09696_ channels.freq1\[9\] _02075_ _02077_ _02078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xrebuffer30 _04162_ net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer41 _06896_ net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_68_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08647_ _01134_ _00040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10289__I _02371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14984__I _06952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08578_ net17 _01093_ _01094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_176_3650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_137_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_137_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10540_ _02798_ _02753_ _02799_ _02800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15536__A1 channels.sample2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_172_3569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10471_ _02695_ _02730_ _02731_ _02732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_157_Right_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_162_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12210_ _04215_ _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_121_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13190_ _05193_ _05194_ _05195_ _05196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12141_ _04152_ _00520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12072_ channels.env_counter\[0\]\[5\] _04114_ _04116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_38_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15900_ _07781_ _07782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_159_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11023_ _03246_ _03247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_99_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16880_ _00949_ _00964_ _00965_ _00966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_15831_ spi_dac_i.counter\[0\] _07717_ _07718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_12974_ _04976_ _04977_ _04980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_63_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15762_ _07332_ _07671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__16595__B _08313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17501_ _00571_ clknet_leaf_14_clk filters.high\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14713_ _06706_ _06691_ _06707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_11925_ _04007_ _04008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14027__A1 _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15693_ _07450_ _07620_ _07621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_169_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09129__S1 _01304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17432_ _00502_ clknet_leaf_182_clk channels.accum\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14644_ _06560_ _06637_ _06638_ _06639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11856_ _03945_ _03946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__15775__A1 _07295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10807_ _03059_ _03060_ _03061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17363_ _00433_ clknet_leaf_97_clk channels.pw2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14575_ _06569_ _06570_ _06571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_60_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09454__A1 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11787_ _03846_ _03851_ _03877_ _03836_ _03878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_83_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16314_ _08154_ _00691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_82_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10738_ _02638_ _02994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13526_ _05531_ _05432_ _05532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_137_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17294_ _00364_ clknet_leaf_187_clk channels.accum\[1\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16245_ _07923_ _08114_ _00662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_24_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13457_ _05327_ _05328_ _05463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_36_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10669_ _02895_ _02926_ _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_113_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_124_Right_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_97_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12408_ _04339_ net34 _04414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_97_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16176_ _08049_ _08050_ _08051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13388_ _05392_ _04933_ _05393_ _05394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_11_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12761__A1 _04714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12339_ _04343_ _04344_ _04345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_15127_ _07090_ _07091_ _07092_ _07093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_11_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_58_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15058_ _07010_ _07025_ _07027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__15674__B filters.sample_buff\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14009_ _06007_ _06009_ _06010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_177_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09550_ _01904_ _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08501_ _01029_ _00132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_144_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10827__A1 _01977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09481_ channels.atk_dec3\[0\] _01867_ _01869_ channels.sus_rel2\[0\] _01871_ channels.freq3\[0\]
+ _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__09693__A1 channels.freq1\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14018__A1 _06014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10055__A2 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_115_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_132_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09817_ _02162_ _02164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_5_10__f_clk clknet_3_2_0_clk clknet_5_10__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__12499__I _04406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14257__A1 _05982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09748_ _01777_ _02107_ _02115_ _00164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_69_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09679_ channels.freq2\[15\] _01997_ _01887_ channels.freq1\[15\] _02063_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_69_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09684__A1 filters.res_filt\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13480__A2 _05208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11710_ _03797_ _03799_ _03800_ _03791_ _03801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_97_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11491__A1 _03513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_174_3609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12690_ _04695_ _04696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_167_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09601__I _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11641_ _03734_ _03735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_83_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13232__A2 _05237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14360_ _06354_ _06355_ _06357_ _06358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_181_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11572_ _03666_ _03680_ _03686_ _00417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_119_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_119_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_135_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13311_ _05314_ _05315_ _05316_ _05317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_10523_ _01089_ _02784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14291_ _06288_ _06183_ _06289_ _06290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_107_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16030_ _07909_ _07818_ _07910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_13242_ _04255_ _04864_ _04491_ _04471_ _05248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10454_ _02685_ _02710_ _02600_ _02714_ _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__14732__A2 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13173_ _03186_ _05179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_10385_ _02644_ _02645_ _02646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12124_ channels.accum\[3\]\[10\] _04144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12055_ _04103_ _04104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16932_ _00011_ clknet_leaf_193_clk channels.ring_outs\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_53_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11006_ _03230_ _03231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_16863_ _03746_ _00941_ _00950_ _00951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_15814_ _06879_ _07698_ _07708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12202__I _04207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16794_ _00899_ _00896_ _00900_ _00901_ _00817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_73_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15745_ _06401_ _07652_ _07659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12957_ _04769_ _04962_ _04763_ _04963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_172_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11908_ _03891_ _03892_ _03899_ _03991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11482__A1 _02289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15676_ _07600_ _07605_ _07606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_23_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12888_ _04893_ _04469_ _04696_ _04378_ _04894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_17415_ _00485_ clknet_leaf_134_clk channels.env_counter\[0\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14627_ _06620_ _06621_ _06622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11839_ _03902_ _03903_ _03930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_23_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17346_ _00416_ clknet_leaf_98_clk channels.freq3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14558_ _05510_ _06005_ _06554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14971__A2 channels.sample3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13509_ _04705_ _05074_ _05515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17277_ _00347_ clknet_leaf_169_clk channels.accum\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14489_ _06480_ _06483_ _06485_ _06486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_113_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16228_ _08088_ _08091_ _08100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_77_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16159_ _07983_ _08008_ _08009_ _07879_ _08025_ _08034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_11_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08981_ _01442_ _01443_ _01444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09038__S0 _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14239__A1 _04504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09602_ filters.cutoff_lut\[13\] _01988_ _01989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09533_ _01875_ _01920_ _01921_ _01922_ _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_108_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09666__A1 filters.hp vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11951__I _04011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09210__S0 _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09666__B2 channels.sus_rel1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09464_ _01789_ _01853_ _01854_ _01855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__15739__A1 _07653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17237__CLK clknet_5_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09421__I _01813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_164_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09395_ _01792_ _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_163_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09969__A2 _02265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12725__A1 _04728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10200__A2 _02455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10170_ channels.pw1\[7\] _02430_ _02431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__14478__A1 _05982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_167_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08500__I _01024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13860_ _05547_ _05862_ _05863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_96_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_159_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12811_ _04816_ _04817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09657__A1 channels.ctrl_reg2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13791_ _04525_ _05793_ _05794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09657__B2 channels.atk_dec2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15530_ filters.sample_buff\[1\] _07461_ _07451_ _07470_ _07471_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_12742_ _04719_ _04746_ _04747_ _04748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_69_Right_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11082__B _03302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09409__A1 filters.lp vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15461_ _07395_ _07399_ _07406_ _07407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_12673_ _04608_ _04609_ _04679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_190_clk clknet_5_22__leaf_clk clknet_leaf_190_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08880__A2 _01342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17200_ _00270_ clknet_leaf_168_clk channels.sync_outs\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14412_ _06407_ _06408_ _06409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11216__A1 filters.high\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11624_ _03721_ _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_182_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15489__B _06952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15392_ filters.low\[22\] _06754_ _07344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_108_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17131_ _00201_ clknet_leaf_127_clk channels.ctrl_reg2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_167_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12964__A1 _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11555_ _01812_ _03675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_14343_ _06339_ _06340_ _06341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_80_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10506_ _02765_ _02766_ _02767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_14274_ _06257_ _06272_ _06273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_17062_ _00132_ clknet_leaf_177_clk filters.res_filt\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_94_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11486_ channels.freq1\[0\] _03626_ _03627_ _03628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12716__A1 _03288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16013_ _07777_ _07890_ _07767_ _07893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_122_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13225_ _04385_ _05231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10437_ _02684_ _02514_ _02607_ _02698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_55_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_78_Right_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13156_ _05160_ _05161_ _05162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_0_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10368_ _02598_ _02628_ _02601_ _02629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_27_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12107_ _04135_ _00503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_104_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13087_ _04764_ _05092_ _05093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10299_ _01328_ _02559_ _02560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12038_ channels.env_counter\[1\]\[11\] _04091_ _04095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16915_ _00957_ channels.exp_periods\[0\]\[0\] _00987_ _00988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_16846_ tt_um_rejunity_sn76489.clk_counter\[3\] _00932_ _00935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16777_ _02272_ _00889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09648__A1 _02030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13989_ _05989_ _05990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_87_Right_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_125_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15728_ _03282_ _07643_ _07644_ _07647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_158_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15659_ channels.sample2\[11\] _03225_ _07589_ _03234_ _07590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_173_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_181_clk clknet_5_19__leaf_clk clknet_leaf_181_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_91_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09180_ channels.lfsr\[3\]\[4\] _01624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_69_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14944__A2 _06910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17329_ _00399_ clknet_leaf_87_clk channels.pw1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_32_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09820__A1 channels.freq2\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_96_Right_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16802__I _00905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_149_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08964_ channels.accum\[0\]\[9\] channels.accum\[1\]\[9\] channels.accum\[2\]\[9\]
+ channels.accum\[3\]\[9\] _01148_ _01163_ _01428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_45_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08895_ _01354_ _01355_ _01363_ _01364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09887__A1 channels.atk_dec2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input17_I rst vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_3_Left_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13435__A2 _05281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12238__A3 _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09639__B2 channels.ctrl_reg3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09516_ _01894_ _01897_ _01902_ _01906_ _01907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_78_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09447_ _01837_ _01838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_109_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_172_clk clknet_5_24__leaf_clk clknet_leaf_172_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_148_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09378_ filters.res_filt\[3\] _01749_ _01763_ _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11340_ _03533_ _03534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_61_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_105_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_169_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11271_ _03465_ _03480_ _03481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__16712__I _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15360__A2 _06599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13010_ _04993_ _05015_ _05016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_162_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10222_ _02432_ _02453_ _02475_ _02482_ _02483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_24_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10185__A1 channels.pw1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_8__f_clk clknet_3_2_0_clk clknet_5_8__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11856__I _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10153_ _02404_ _02409_ _02413_ _01553_ _02414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_33_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09326__I _01728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10084_ clk_trg\[0\] _02350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_50_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14961_ _06918_ _06933_ _00559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16700_ _08419_ _08439_ _00792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13912_ _04451_ _04862_ _05914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17680_ _00750_ clknet_leaf_69_clk tt_um_rejunity_sn76489.tone\[1\].gen.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11685__A1 _03535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14892_ _06868_ _06870_ _00553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_96_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16631_ _01689_ _08386_ _08387_ _01691_ _00775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_13843_ _05762_ _05765_ _05845_ _05846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XTAP_TAPCELL_ROW_18_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14623__A1 _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13426__A2 _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16562_ _08336_ _08341_ _08342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_97_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13774_ _05689_ _05691_ _05776_ _05777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10986_ filters.high\[0\] _03210_ _03211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09061__I _01257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15513_ _03263_ _07453_ _07454_ _03219_ _07455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_12725_ _04728_ _04259_ _04695_ _04729_ _04731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_16493_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[3\] _08268_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[3\]
+ _08284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_48_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_163_clk clknet_5_28__leaf_clk clknet_leaf_163_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_155_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10000__I _02290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15444_ _07386_ _07390_ _07392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_84_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10660__A2 _02872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12656_ _04652_ _04660_ _04661_ _04662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_127_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12937__A1 _04863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11607_ _03677_ _03703_ _03709_ _00429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_53_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10935__I _01320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12587_ _03272_ _04242_ _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15375_ filters.low\[20\] _06599_ _07328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09802__A1 channels.sus_rel1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17114_ _00184_ clknet_leaf_116_clk channels.sus_rel1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__16679__A2 _08244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14326_ _06322_ _06323_ _06324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_11538_ channels.freq2\[1\] _03659_ _03660_ _03663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_123_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14851__B _06717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17045_ _00115_ clknet_leaf_238_clk channels.lfsr\[1\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14257_ _05982_ _06086_ _06098_ _06256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11469_ _03618_ _03615_ _01539_ _03616_ _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13362__A1 _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12165__A2 _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13208_ _03270_ _04240_ _05106_ _05214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_1_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14188_ _03330_ _06080_ _06185_ _06187_ _00532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13139_ _05107_ _05145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__15103__A2 _01927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input9_I bus_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09869__A1 _02131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13981__I _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12468__A3 _04390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11676__A1 _01168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08680_ _01163_ _01164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_174_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16829_ _03496_ _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_152_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_178_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09301_ _01726_ _01727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_85_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16367__A1 channels.ch3_env\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_154_clk clknet_5_29__leaf_clk clknet_leaf_154_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_159_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09232_ _01664_ _01659_ _01668_ _01651_ _00091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_111_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10651__A2 _02622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09163_ channels.lfsr\[2\]\[3\] _01609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_161_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_10__f_clk_I clknet_3_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11600__A1 channels.pw3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09094_ channels.accum\[0\]\[20\] _01547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__15857__B _07740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14761__B _06734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13353__A1 _04500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09557__B1 _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10580__I _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09996_ channels.ctrl_reg3\[7\] _02283_ _02284_ _02288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_181_3741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08947_ channels.freq3\[8\] _01397_ _01412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14853__B2 _06752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11667__A1 channels.sus_rel1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08878_ _01336_ _01262_ _01348_ _01318_ _00057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_4_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11625__B _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14605__A1 _03396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10840_ _03092_ _03093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_67_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10771_ _02993_ _02997_ _03026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xclkbuf_leaf_145_clk clknet_5_30__leaf_clk clknet_leaf_145_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_55_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12510_ _04497_ _04502_ _04515_ _04516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_13490_ _05495_ _05345_ _05496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_164_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12441_ _04446_ _04447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_164_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13592__A1 _04220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12372_ _04377_ _04378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15160_ _07101_ _07123_ _07124_ _07125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11323_ _03519_ _03520_ _03521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_16_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14111_ _03413_ _04488_ net58 _06111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_26_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15091_ _07056_ _07024_ _07058_ _07059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__16442__I _08242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16530__A1 _08242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11254_ _03454_ _03463_ _03464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_120_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14042_ _05914_ _05915_ _06043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10205_ _02427_ channels.pw2\[1\] _02465_ _01096_ _02466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_63_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11185_ _03335_ _03400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10136_ _01071_ _02397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15993_ _07839_ _07833_ _07865_ _07873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_66_Left_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_89_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17732_ _00802_ clknet_leaf_64_clk tt_um_rejunity_sn76489.control_tone_freq\[1\]\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10067_ filters.cutoff_lut\[12\] _02332_ _02335_ _02339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14944_ _04214_ _06910_ _06914_ _06916_ _06917_ _00558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_17663_ _00733_ clknet_leaf_57_clk tt_um_rejunity_sn76489.noise\[0\].gen.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14875_ _06840_ _06847_ _06855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10330__A1 _02522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16614_ _08377_ _08382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12210__I _04215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13826_ _04445_ _05828_ _05829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17594_ _00664_ clknet_leaf_39_clk spi_dac_i.spi_dat_buff_0\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10881__A2 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16545_ _08322_ _08327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_156_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_136_clk clknet_5_31__leaf_clk clknet_leaf_136_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_134_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13757_ _03269_ _05545_ _05760_ _05653_ _00528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_10969_ _03193_ _03194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_128_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12708_ _04186_ _04713_ _04714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_100_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16476_ _08268_ _08269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_17_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13688_ _05689_ _05691_ _05692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_72_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_75_Left_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_80_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15427_ _07375_ _07376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_31_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12639_ _04644_ _04645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_143_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15358_ _07030_ _07312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08685__S1 _01168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14309_ _06253_ _06273_ _06307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15324__A2 _07062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15289_ _05852_ _07233_ _07248_ _07249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_17028_ _00005_ clknet_leaf_240_clk filters.res_lut\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_146_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09850_ _01765_ _02187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__15088__A1 _04992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_84_Left_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08801_ _01273_ _01274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11361__A3 _03531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09781_ _02137_ _02138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08732_ _01184_ _01190_ _01215_ _01216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_1_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08663_ _01146_ _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_178_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16588__A1 _08333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_120_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08594_ channels.lfsr\[3\]\[1\] _01108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10872__A2 _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_209_clk_I clknet_5_17__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14063__A2 _05967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_127_clk clknet_5_27__leaf_clk clknet_leaf_127_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__16527__I _01822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_138_Right_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_113_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_93_Left_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_174_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09215_ channels.lfsr\[1\]\[9\] _01654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16760__A1 _08456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09146_ channels.lfsr\[2\]\[1\] _01594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_118_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09077_ channels.accum\[0\]\[18\] _01532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_102_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_135_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_9_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09979_ channels.ctrl_reg3\[0\] _02276_ _02277_ _02278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10560__A1 _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12990_ _04994_ _04995_ _04996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08505__A1 _01008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09604__I _01866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11941_ channels.env_counter\[2\]\[2\] _04013_ _04022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_170_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12030__I _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14660_ _06540_ _06559_ _06654_ _06655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11872_ _03939_ _03958_ _03959_ _00444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_1265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13611_ _05607_ _05615_ _05616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10823_ _03074_ _03076_ _03077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_95_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_118_clk clknet_5_26__leaf_clk clknet_leaf_118_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_14591_ _06584_ _06585_ _06586_ _06587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_45_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_105_Right_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13801__A2 _05260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16330_ _03958_ _08158_ _08164_ _00697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13542_ _05546_ _05547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10754_ _03008_ _03009_ _03010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16261_ filters.sample_buff\[8\] _08125_ _08122_ spi_dac_i.spi_dat_buff_0\[4\] spi_dac_i.spi_dat_buff_0\[5\]
+ _08119_ _08126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_82_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13473_ _03350_ _04192_ _05220_ _05479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_10685_ _02938_ _02941_ _02942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_153_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15212_ _03394_ _07162_ _07175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_164_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12424_ _04362_ _04428_ _04430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16192_ _07882_ _07887_ _08066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_124_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15143_ _07107_ _07108_ _07109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_23_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12355_ _04352_ _04359_ _04361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11306_ _03507_ _03508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12286_ _04291_ _04292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15074_ _07019_ _07020_ _07042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__13868__A2 _05643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11237_ _03447_ _03448_ _03449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14025_ _05927_ _05932_ _06025_ _06026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12540__A2 _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11168_ _03374_ _03378_ _03383_ _03230_ _03384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__10551__A1 _02544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10119_ channels.ctrl_reg1\[5\] _01286_ _02380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_15976_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[0\] _07765_ _07857_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_141_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11099_ filters.high\[5\] _03210_ _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17715_ _00785_ clknet_leaf_68_clk tt_um_rejunity_sn76489.tone\[0\].gen.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_175_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14927_ _06720_ _06893_ _06902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16775__C _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17646_ _00716_ clknet_leaf_51_clk tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_180_clk_I clknet_5_19__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10854__A2 _03104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14858_ _06836_ _06839_ _06840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_82_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13809_ _05719_ _05737_ _05812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_109_clk clknet_5_15__leaf_clk clknet_leaf_109_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_17577_ _00647_ clknet_leaf_33_clk spi_dac_i.counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_60_clk_I clknet_5_8__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14789_ _06689_ _06777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_58_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16528_ _08310_ _08312_ _08313_ _00746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_128_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_195_clk_I clknet_5_23__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16459_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[5\] _08251_ _08255_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_143_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09000_ channels.accum\[0\]\[11\] _01461_ _01462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12359__A2 _04327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_7_0_clk clknet_0_clk clknet_3_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_182_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_75_clk_I clknet_5_14__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13020__A3 _05000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_170_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09902_ channels.atk_dec2\[6\] _02220_ _02217_ _02223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_113_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_130_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_133_clk_I clknet_5_31__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09833_ _01750_ _02174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09764_ channels.atk_dec1\[0\] _02126_ _02120_ _02127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_13_clk_I clknet_5_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09424__I net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08715_ _01198_ _01199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_154_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09695_ _01808_ _02077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xrebuffer20 _05151_ net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_96_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_148_clk_I clknet_5_31__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer31 _04177_ net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_96_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xrebuffer42 _04493_ net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08646_ channels.env_vol\[3\]\[4\] _01134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15233__A1 _03410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12785__I _04783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08577_ _01068_ _01093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA__15784__A2 _07682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_176_3651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14992__B1 channels.sample2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_137_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15536__A2 _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10470_ _02652_ _02673_ _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_40_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09129_ channels.lfsr\[0\]\[22\] channels.lfsr\[1\]\[22\] channels.lfsr\[2\]\[22\]
+ channels.lfsr\[3\]\[22\] _01201_ _01304_ _01578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_32_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16921__S _00987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08974__A1 _01427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12140_ channels.accum\[3\]\[18\] _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_60_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12071_ _04029_ _04113_ _04115_ _00487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11022_ filters.filter_step\[2\] _03246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__16249__C2 _07728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15830_ spi_dac_i.counter\[4\] spi_dac_i.counter\[3\] _07717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_99_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15761_ _07639_ _07670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_12973_ _04957_ _04956_ _04958_ _04979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_17500_ _00570_ clknet_leaf_249_clk filters.high\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14712_ _06700_ _06706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_11924_ _04006_ _04007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10836__A2 _02840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15692_ _07616_ _07613_ _07618_ _07620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_87_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17431_ _00501_ clknet_leaf_153_clk channels.adsr_state\[1\]\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14643_ _06563_ _06591_ _06638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11855_ _03778_ _03934_ _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15775__A2 _07631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14822__I1 filters.band\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12589__A2 _04171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10806_ _03037_ _03041_ _03060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17362_ _00432_ clknet_leaf_93_clk channels.pw2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_14574_ _04893_ _05687_ _06570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11786_ _03803_ _03858_ _03868_ _03877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09454__A2 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16313_ channels.env_counter\[3\]\[12\] _08154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_165_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13525_ _05527_ _05530_ _05531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10737_ _02602_ _02776_ _02993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17293_ _00363_ clknet_leaf_188_clk channels.accum\[2\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_137_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13538__A1 _03730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16244_ filters.sample_buff\[3\] _07722_ _07728_ spi_dac_i.spi_dat_buff_0\[0\] _08114_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_67_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13456_ _05327_ _05328_ _05462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_82_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_149_Left_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10668_ _02914_ _02925_ _02926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_24_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12407_ _04381_ _04410_ _04412_ _04413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XTAP_TAPCELL_ROW_97_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16175_ _07909_ _07820_ _07823_ _07847_ _07908_ _08050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_141_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13387_ _04877_ _04907_ _05393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_11_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10599_ _02856_ _02857_ _02858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08965__A1 _01427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15126_ _07079_ _07081_ _07092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12338_ _03316_ _04164_ _04199_ _04344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_58_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15057_ _07010_ _07025_ _07026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_12269_ _04274_ _04187_ _04275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_75_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14008_ _04487_ _06008_ _06009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10524__A1 channels.sample3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_158_Left_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_170_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09244__I _01604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15959_ _07839_ _07833_ _07840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12816__A3 _04444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08500_ _01024_ _01029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09480_ _01870_ _01871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_114_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17629_ _00699_ clknet_leaf_210_clk channels.env_vol\[1\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15766__A2 _07670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_154_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_154_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_167_Left_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_160_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_156_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13529__A1 _05534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17016__CLK clknet_5_16__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_171_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_115_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12201__A1 filters.res_lut\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09816_ _02162_ _02163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_119_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16696__B _01823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09747_ channels.ctrl_reg1\[3\] _02108_ _02113_ _02115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09678_ filters.mode_vol\[7\] _02014_ _02001_ channels.freq2\[7\] _02062_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_119_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15206__A1 _07146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08629_ _01125_ _00031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_96_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15757__A2 _07632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11640_ _03733_ _03734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_92_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11571_ channels.freq3\[3\] _03681_ _03682_ _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_181_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13310_ _04477_ _04781_ _04784_ _04267_ _05316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_10522_ _02733_ _02736_ _02782_ _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_52_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14290_ _06287_ _06179_ _06289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_150_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13241_ _05200_ _05245_ _05246_ _05247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10453_ _02704_ _02706_ _02711_ _02713_ _02714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_21_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10384_ _02590_ _02645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13172_ _05173_ _05177_ _05178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__15775__B _07648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12123_ _04143_ _00511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_62_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16931_ _01766_ _00923_ _00996_ _00919_ _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_12054_ _03744_ _04005_ _04103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_53_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11005_ _03229_ _03230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_99_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16862_ _03745_ _03752_ _03775_ _00950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__15445__A1 _06909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09064__I _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15813_ _07706_ _07707_ _00637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_70_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16793_ _02102_ _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_88_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10003__I _02293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15744_ _07655_ _07658_ _00617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12956_ _04208_ _04766_ _04962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_133_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11907_ _03844_ _03867_ _03875_ _03990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11482__A2 _01954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15675_ _07603_ _07604_ _07605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_34_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10938__I _01460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12887_ _04316_ _04893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_17414_ _00484_ clknet_leaf_132_clk channels.env_counter\[0\]\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14626_ _06565_ _06573_ _06621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11838_ _01584_ _03921_ _03922_ _03928_ _03929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_8_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17345_ _00415_ clknet_leaf_96_clk channels.freq3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_16_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14557_ _05512_ _05796_ _06553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11769_ _03850_ _03859_ _03860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_138_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_40_clk clknet_5_3__leaf_clk clknet_leaf_40_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_71_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13508_ _05342_ _05511_ _05513_ _05514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_67_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17276_ _00346_ clknet_leaf_181_clk channels.accum\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14488_ _06484_ _05560_ _06485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16227_ _08097_ _08099_ _00659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_126_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13439_ _04561_ _05370_ _05445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16158_ _08007_ _08031_ _08032_ _08033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_51_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10745__A1 _02657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15109_ _07073_ _07074_ _07075_ _07076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_110_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16089_ _07964_ _07936_ _07966_ _07967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08980_ channels.accum\[0\]\[10\] channels.accum\[1\]\[10\] channels.accum\[2\]\[10\]
+ channels.accum\[3\]\[10\] _01149_ _01164_ _01443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XTAP_TAPCELL_ROW_110_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09038__S1 _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09363__A1 _01757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09601_ _01956_ _01988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09532_ channels.pw1\[1\] _01885_ _01887_ channels.freq1\[9\] _01922_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13998__A1 _05905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_108_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09210__S1 _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09463_ _00997_ _01784_ _01854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_94_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13224__I _04784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09394_ _01792_ _01793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_172_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14175__A1 _05877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12725__A2 _04259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10200__A3 channels.pw3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_98_clk clknet_5_13__leaf_clk clknet_leaf_98_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_100_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12810_ filters.cutoff_lut\[14\] _04441_ _04816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_13790_ _05690_ _05793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09612__I _01881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12741_ _04727_ _04745_ _04747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_96_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16927__A1 _01741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15460_ _07383_ _06767_ _07396_ _07406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_38_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12672_ _04674_ _04675_ _04677_ _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_38_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14402__A2 _06399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14411_ _06372_ _06387_ _06408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11623_ _02100_ _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_33_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15391_ _07327_ _06716_ _07343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_22_clk clknet_5_3__leaf_clk clknet_leaf_22_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_17130_ _00200_ clknet_leaf_117_clk channels.ctrl_reg2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_64_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12964__A2 _04966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14342_ _04318_ _05500_ _06340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11554_ _03673_ _03669_ _03674_ _00411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_167_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_135_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_1307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10505_ _02662_ _02623_ _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17061_ _00131_ clknet_leaf_176_clk filters.res_filt\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14273_ _06270_ _06271_ _06272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11485_ _03516_ _03627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_123_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16012_ _07769_ _07857_ _07892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_150_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13224_ _04784_ _05230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12716__A2 _04316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10436_ _02684_ _02628_ _02686_ _02697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_100_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_55_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09593__A1 channels.pw2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09593__B2 channels.atk_dec1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13155_ _03363_ _04315_ _04271_ _05161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10367_ _02528_ _02628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_104_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12106_ channels.accum\[3\]\[1\] _04135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13086_ _05091_ _05092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10298_ channels.env_vol\[0\]\[1\] channels.env_vol\[1\]\[1\] _01144_ _02559_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_89_clk clknet_5_12__leaf_clk clknet_leaf_89_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12037_ _04056_ _04090_ _04094_ _00474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12213__I _04218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16914_ _00986_ _00987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_18_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16845_ tt_um_rejunity_sn76489.clk_counter\[3\] _00932_ _00934_ _00835_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__16091__A1 _07956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16776_ net9 _00886_ _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13988_ _05796_ _05989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_158_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15727_ _05862_ _07637_ _07646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_158_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11455__A2 _03605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12939_ _04858_ _04945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15658_ _03421_ _07563_ _07588_ _03224_ _07589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_133_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14609_ _06499_ _06501_ _06605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15589_ channels.sample3\[6\] _07513_ _07525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_13_clk clknet_5_6__leaf_clk clknet_leaf_13_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_172_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17328_ _00398_ clknet_leaf_87_clk channels.pw1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_16_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_32_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17259_ _00329_ clknet_leaf_72_clk tt_um_rejunity_sn76489.control_tone_freq\[0\]\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_149_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_149_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15657__A1 _02056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08963_ _01424_ _01426_ _01427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_80_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15862__C _07710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08894_ _01350_ _01347_ _01356_ _01363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_127_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_127_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12891__A1 _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15434__I _01932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09432__I _01822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09639__A2 _01937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13435__A3 _05372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09515_ channels.sample3\[4\] _01904_ _01905_ clk_trg\[0\] _01906_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_116_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12643__B2 _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09446_ _01836_ _01828_ _01832_ _01837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_140_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09377_ _01776_ _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14148__A1 _06015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15896__A1 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[0\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11270_ _03466_ _03479_ _03480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_160_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_104_Left_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10221_ _02476_ _02477_ _02451_ _02481_ _02482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__15648__A1 filters.sample_buff\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10152_ _02410_ _02411_ _02412_ _02413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10083_ _01933_ _02349_ _00265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_50_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14960_ filters.high\[1\] _06919_ _06930_ _06932_ _06933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_50_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13911_ _04324_ _05078_ _05913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__11685__A2 _03771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14891_ _06520_ _06869_ _06860_ _06870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16630_ _01681_ _08386_ _08387_ _01684_ _00774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_13842_ _05782_ _05785_ _05844_ _05845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_96_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_113_Left_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_18_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16561_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[3\] _08327_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[3\]
+ _08341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13773_ _04597_ _05775_ _05692_ _05776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_168_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10985_ _03209_ _03210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_139_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15512_ channels.sample3\[0\] _07453_ _07454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12724_ _04728_ _04695_ _04729_ _04259_ _04730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_16492_ _08279_ _08283_ _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_139_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15443_ _07386_ _07390_ _07391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12655_ _04623_ _04624_ _04612_ _04661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_154_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11606_ channels.pw3\[7\] _03704_ _03705_ _03709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15374_ filters.low\[21\] _07327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12586_ _04581_ _04582_ _04592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_4_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10948__A1 channels.sample1\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17113_ _00183_ clknet_leaf_116_clk channels.sus_rel1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14325_ _04820_ _04924_ _06323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11537_ _01755_ _03662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_128_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17044_ _00114_ clknet_leaf_228_clk channels.lfsr\[1\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09015__B1 _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14256_ _06254_ _06096_ _06095_ _06255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_151_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11468_ channels.accum\[1\]\[18\] _03618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09566__A1 channels.ch3_env\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13207_ _03285_ _04195_ _04880_ _05213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09566__B2 channels.freq1\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10419_ _02607_ _02645_ _02680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14187_ _06186_ _06187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11399_ channels.accum\[2\]\[14\] _03577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10176__A2 channels.pw2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09517__I _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11268__B _03236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13138_ _04368_ _04881_ _05144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09318__A1 _01657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14311__A1 _06197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13069_ _05074_ _05075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_2_clk clknet_5_1__leaf_clk clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_144_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_119_Right_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_144_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12873__A1 filters.cutoff_lut\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16064__A1 _07929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16828_ _00923_ _00924_ _01823_ _00828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_75_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16759_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[7\] _00873_ _00871_ _00875_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_85_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_122_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09300_ _01725_ _01726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_174_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09231_ _01665_ _01666_ _01658_ _01667_ _01305_ _01656_ _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_150_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09162_ _01600_ _01592_ _01608_ _01599_ _00081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_17_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10939__A1 channels.sample1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09093_ _01540_ _01545_ _01546_ _00074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09557__A1 channels.sus_rel1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09557__B2 channels.sample3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13353__A2 _05092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09427__I _01818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09995_ _02240_ _02282_ _02287_ _00239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_177_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08946_ _01410_ _01411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_181_3742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08877_ _01337_ _01344_ _01347_ _01348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_4_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16055__A1 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[2\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14605__A2 _06067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12616__A1 _04541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10770_ _03023_ _03024_ _03025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09429_ _01819_ _01802_ _01820_ _00140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_35_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12919__A2 _04924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12440_ _04445_ _04446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13041__A1 _04952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09796__A1 channels.sus_rel1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13592__A2 _04926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12371_ _04376_ _04377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14110_ _03397_ _04402_ _05106_ _06110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11322_ _01811_ _03495_ _03520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_132_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15090_ _07057_ _07058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_50_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15339__I filters.low\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14041_ _06026_ _06041_ _06042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_11253_ _03461_ _03463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10204_ _01072_ channels.pw1\[1\] _02465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_30_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11184_ _03394_ _03395_ _03398_ _03232_ _03399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_101_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10135_ _02391_ _02392_ _02396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_15992_ _07838_ _07866_ _07872_ _00651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_89_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_89_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17731_ _00801_ clknet_leaf_63_clk tt_um_rejunity_sn76489.control_tone_freq\[1\]\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10066_ _02316_ _02331_ _02338_ _00259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14943_ _02353_ _06917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_121_Left_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17662_ _00732_ clknet_leaf_58_clk tt_um_rejunity_sn76489.noise\[0\].gen.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14874_ _06852_ _06853_ _06854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_89_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10330__A2 _02590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09072__I _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13825_ _05469_ _05828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16613_ _08380_ _08381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17593_ _00663_ clknet_leaf_38_clk spi_dac_i.spi_dat_buff_0\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12607__A1 _03256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15802__I _07355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16544_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[1\] _08326_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13756_ _05547_ _05759_ _05760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_174_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16349__A2 _01317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10968_ _03192_ _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_128_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12707_ _04712_ _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_73_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_100_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16475_ _08260_ _08268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_63_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13687_ _04400_ _05690_ _05691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10633__A3 _02890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10899_ channels.sample2\[2\] _03143_ _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15426_ _07372_ _06852_ _07375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_130_Left_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12638_ _04643_ _04644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_80_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15357_ _07035_ _07309_ _07311_ _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_5_2__f_clk_I clknet_3_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16633__I _08382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12569_ _04231_ _04575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_81_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_170_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11594__A1 _03664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10397__A2 _02657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14308_ _06194_ _06252_ _06306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15288_ _07247_ _07248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__16521__A2 _08282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17027_ _00004_ clknet_leaf_240_clk filters.res_lut\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14239_ _04504_ _05989_ _06238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_146_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08800_ _01248_ _01272_ _01273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_42_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09780_ _01751_ _02137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11361__A4 _03549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08731_ _01197_ _01212_ _01214_ _01215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_147_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09711__A1 channels.freq1\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08662_ _01145_ _01146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_178_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_120_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08593_ _01107_ _00013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_163_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_120_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13271__A1 _05184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10085__A1 _02088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09214_ channels.lfsr\[0\]\[9\] _01653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_157_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09778__A1 channels.atk_dec1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09145_ _01580_ _01589_ _01592_ _01593_ _00079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_133_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_135_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09076_ _01531_ _00072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_135_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09157__I _01201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09978_ _02254_ _02277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_157_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08929_ _01383_ _01262_ _01395_ _01318_ _00061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12837__A1 _04732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16919__S _00987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08505__A2 _01019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11940_ _04019_ _04020_ _04021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12311__I _04316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_169_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11871_ channels.env_vol\[0\]\[3\] _03942_ _03959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16718__I _08445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13610_ _05610_ _05614_ _05615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__15251__A2 channels.sample1\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10822_ _03075_ _03044_ _03076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_14590_ _05624_ _05091_ _06586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09620__I _01844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10076__A1 filters.cutoff_lut\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11273__B1 _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13541_ _05543_ _05546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10753_ _02986_ _03007_ _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16260_ _07741_ _08125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13472_ _04511_ _04445_ _05478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10684_ _02839_ _02919_ _02940_ _02941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_152_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15211_ _03394_ _07162_ _07174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09769__A1 channels.atk_dec1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12423_ _04362_ _04428_ _04429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_16191_ _07933_ _07891_ _07932_ _08065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_164_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15142_ _01746_ channels.sample1\[7\] _07108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12354_ _04352_ _04359_ _04360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11305_ _01812_ _03491_ _03492_ _03495_ _03507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_132_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13317__A2 _05237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15073_ _07019_ _07020_ _07041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_12285_ _04290_ _04291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_65_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11328__A1 _02103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14024_ _05922_ _05926_ _06025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_31_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11236_ _03436_ _03438_ _03448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11167_ _03382_ _03383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_101_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10118_ _01527_ _02378_ _02379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__12828__A1 _04324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15975_ _07767_ _07770_ _07856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_141_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11098_ _03310_ _03217_ _03317_ _03228_ _03318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_141_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17714_ _00784_ clknet_leaf_67_clk tt_um_rejunity_sn76489.tone\[0\].gen.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10049_ _01813_ _02326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_14926_ _06720_ _06893_ _06901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_175_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11500__A1 _02324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17645_ _00715_ clknet_leaf_49_clk tt_um_rejunity_sn76489.chan\[3\].attenuation.in
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14857_ _06837_ _03474_ _06838_ _06839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_26_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13253__S _03185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13808_ _05789_ _05810_ _05811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_17576_ _00646_ clknet_leaf_33_clk spi_dac_i.counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14788_ _06761_ _06774_ _06776_ _00543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10067__A1 filters.cutoff_lut\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16527_ _01822_ _08313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_129_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13739_ _05660_ _05742_ _05743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_46_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16458_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[5\] _08251_ _08254_ _00735_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_144_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15409_ _07336_ _07345_ _07353_ _07359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_16389_ _08202_ _08203_ _08200_ _00717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11567__A1 channels.freq3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_130_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13308__A2 _04800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09901_ _02155_ _02219_ _02222_ _00210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_112_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_113_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_113_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_130_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09832_ _02155_ _02170_ _02173_ _00190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09932__A1 channels.sus_rel2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_171_Right_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09763_ _02124_ _02126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08714_ channels.exp_counter\[0\]\[3\] channels.exp_counter\[1\]\[3\] channels.exp_counter\[2\]\[3\]
+ channels.exp_counter\[3\]\[3\] _01178_ _01172_ _01198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_09694_ _01742_ _02074_ _02076_ _00149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13492__A1 _05324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer10 _05431_ net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer21 _04812_ net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_179_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer32 _05411_ net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_83_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_178_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08645_ _01133_ _00039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_178_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_159_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_159_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08576_ channels.clk_div\[0\] _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_178_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_176_3641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_176_3652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09999__A1 _02289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14992__A1 filters.filt_1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14992__B2 filters.filt_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_174_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_40_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09128_ _01573_ _01574_ _01575_ _01576_ _01201_ _01304_ _01577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_161_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12306__I _04311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09059_ _01422_ _01515_ _01516_ _00070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11210__I filters.band\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12070_ channels.env_counter\[0\]\[4\] _04114_ _04115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_240_clk_I clknet_5_18__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16249__A1 filters.sample_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09923__A1 _02234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11021_ _03212_ _03213_ _03243_ _03245_ _03179_ _00307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_TAPCELL_ROW_38_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15472__A2 _06717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15760_ _06728_ _07664_ _07669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12972_ _04976_ _04977_ _04978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10297__A1 _01307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11923_ _02356_ _04005_ _04006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14711_ _06699_ _06606_ _06702_ _06704_ _06705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
X_15691_ _07616_ _07613_ _07618_ _07619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14642_ _06592_ _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_17430_ _00500_ clknet_leaf_159_clk channels.adsr_state\[1\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11854_ _03537_ _03749_ _03944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09350__I _01752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10805_ _03027_ _03036_ _03059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17361_ _00431_ clknet_leaf_97_clk channels.pw2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_14573_ _04452_ _05505_ _06569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11785_ _03863_ _03867_ _03875_ _03876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_138_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_60_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16312_ _08153_ _00690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13524_ _05528_ net44 _05529_ _05530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_10736_ _02954_ _02956_ _02991_ _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_17292_ _00362_ clknet_leaf_155_clk channels.accum\[2\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_16243_ _07924_ _08112_ _08113_ _00661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13455_ _05321_ _05331_ _05460_ _05461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10667_ _02919_ _02924_ _02925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_141_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12406_ _04339_ _04347_ _04411_ _04412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_113_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16174_ _08044_ _08048_ _08049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_97_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13386_ _04877_ _04907_ _05392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_97_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10598_ _02850_ _02855_ _02857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_11_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15125_ _07079_ _07081_ _07091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_142_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12337_ _03383_ _04342_ _04185_ _04343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__12216__I _04221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_58_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15056_ _04992_ _07012_ _07024_ _07025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_103_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12268_ _04273_ _04274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_208_clk_I clknet_5_22__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09914__A1 channels.sus_rel2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14007_ filters.high\[25\] filters.band\[25\] _03187_ _06008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11219_ _03416_ _03432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_12199_ _04183_ _04203_ _04204_ _04205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_37_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15958_ _07807_ _07831_ _07839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13474__A1 _03364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10288__A1 _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14909_ _06719_ _06877_ _06886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_15889_ _07768_ _07769_ _07770_ _07771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17628_ _00698_ clknet_leaf_213_clk channels.env_vol\[1\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17559_ _00629_ clknet_leaf_245_clk filters.low\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_160_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_154_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_154_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10460__A1 _01164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13529__A2 _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_171_3560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13510__I _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_132_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11960__A1 _04019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09905__A1 channels.atk_dec2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09815_ _02123_ _01893_ _02162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09746_ _02112_ _02107_ _02114_ _00163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13465__A1 _04451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10279__A1 _01470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11476__B1 _01568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09677_ channels.freq1\[7\] _02011_ _01936_ channels.sus_rel2\[7\] _02061_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_9_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15206__A2 _07149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08628_ channels.lfsr\[3\]\[18\] _01125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_68_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08559_ _01075_ _01076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14965__A1 _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14944__C _06917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11570_ _03664_ _03680_ _03685_ _00416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_107_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10521_ _02738_ _02781_ _02782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14717__A1 _03422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13240_ _05157_ _05163_ _05246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10452_ _02712_ _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13171_ _05174_ _05175_ _05176_ _05177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__11400__B1 _01503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10383_ _02536_ _02644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13940__A2 _05504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12122_ channels.accum\[3\]\[9\] _04143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16930_ tt_um_rejunity_sn76489.control_noise\[0\]\[2\] _00923_ _00996_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12053_ _04101_ _03732_ _04102_ _00482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_53_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11004_ _03228_ _03229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_53_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16861_ _03768_ _03971_ _00941_ _00948_ _00949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__15791__B _07684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_194_clk_I clknet_5_23__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_70_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15812_ _07395_ _07694_ _07695_ _07707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_70_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16792_ net9 _00897_ _00900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_3_6_0_clk clknet_0_clk clknet_3_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_clkbuf_leaf_74_clk_I clknet_5_9__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12955_ _04956_ _04959_ _04960_ _04961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_73_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15743_ _03345_ _07656_ _07657_ _07658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_137_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11906_ _03860_ _03862_ _03988_ _03989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13208__A1 _03270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15674_ _03450_ _07602_ filters.sample_buff\[12\] _07604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_12886_ _04449_ _04696_ _04378_ _04469_ _04892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__08883__B2 channels.freq1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17413_ _00483_ clknet_leaf_132_clk channels.env_counter\[0\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11837_ _03923_ _03926_ _03927_ _03928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_14625_ _06567_ _06572_ _06620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14956__A1 _05534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_89_clk_I clknet_5_12__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17344_ _00414_ clknet_leaf_100_clk channels.freq3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_126_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14556_ _04575_ _06008_ _06552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11768_ _03837_ _03827_ _03858_ _03859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_132_clk_I clknet_5_31__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08852__C _01303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13507_ _05512_ _05510_ _04758_ _04946_ _05513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_67_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10719_ channels.sample3\[4\] _02975_ _02976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14708__A1 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14487_ filters.band\[27\] _06484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_17275_ _00345_ clknet_leaf_179_clk channels.accum\[2\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11699_ _03788_ _03789_ _03790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_82_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16226_ spi_dac_i.spi_dat_buff_1\[9\] _07924_ _08098_ _08099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13438_ _05335_ _05356_ _05443_ _05444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_153_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xrebuffer1 net43 net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_180_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_248_clk clknet_5_1__leaf_clk clknet_leaf_248_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_16157_ _08026_ _08028_ _08032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_141_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_147_clk_I clknet_5_29__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13369_ _05299_ _05358_ _05374_ _05375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_12_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10745__A2 _02823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15108_ _01746_ channels.sample1\[6\] _07075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16088_ _07896_ _07902_ _07965_ _07966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_11_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_27_clk_I clknet_5_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15039_ _05969_ _06993_ _07008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13695__A1 _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09600_ _01933_ _01987_ _00144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11170__A2 _03385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13447__A1 _05451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09531_ channels.freq2\[1\] _01880_ _01882_ channels.ctrl_reg3\[1\] _01921_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_91_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11458__B1 _01503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13998__A2 _05935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09462_ _01827_ _01853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_78_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_3600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09393_ _01781_ _01791_ _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_171_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10984__A2 _03205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_239_clk clknet_5_16__leaf_clk clknet_leaf_239_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__13922__A2 _05731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09165__I _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16624__A1 _01657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09106__A2 _01556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09729_ _02100_ _02101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_167_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12740_ _04727_ _04745_ _04746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_85_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output23_I net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16927__A2 _00993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12671_ _04676_ _04586_ _04677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_132_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14410_ _06311_ _06371_ _06407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_155_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11622_ _03711_ _03720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_167_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15390_ _07341_ _07342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_108_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14341_ _04378_ _05447_ _06339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11553_ channels.freq2\[5\] _03670_ _03671_ _03674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_37_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10504_ _02643_ _02648_ _02764_ _02765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_17060_ _00130_ clknet_leaf_178_clk filters.res_filt\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_14272_ _06259_ _06269_ _06271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11484_ _03624_ _03626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_162_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16011_ _07890_ _07778_ _07891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12177__A1 _04176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13223_ _04824_ _05229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_123_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13913__A2 _04927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10435_ _02681_ _02682_ _02696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_61_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13154_ _03348_ _04191_ _04375_ _05160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_55_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10366_ _02577_ _02584_ _02627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12105_ _04134_ _00502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_72_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13085_ _04927_ _05091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10297_ _01307_ channels.env_vol\[3\]\[1\] _02557_ _02558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_12036_ channels.env_counter\[1\]\[10\] _04091_ _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16913_ _03744_ _03728_ _01043_ _00986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_18_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10014__I _02290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16844_ tt_um_rejunity_sn76489.clk_counter\[3\] _00932_ _00877_ _00934_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16775_ _07826_ _00885_ _00887_ _02273_ _00812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_13987_ _04630_ _05892_ _05988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14641__A3 _06635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15726_ _07642_ _07645_ _00612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_87_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12938_ _04859_ _04942_ _04943_ _04944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_34_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10663__A1 _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15657_ _02056_ _07563_ _07588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12869_ _04815_ _04839_ _04875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_103_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14608_ _06499_ _06501_ _06604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_50_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15588_ filters.sample_buff\[5\] _07518_ _07524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17327_ _00397_ clknet_leaf_88_clk channels.freq1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14539_ _06415_ _06446_ _06535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17258_ _00328_ clknet_leaf_72_clk tt_um_rejunity_sn76489.control_tone_freq\[0\]\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16209_ _08080_ _08081_ _08082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_70_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17189_ _00259_ clknet_leaf_78_clk filters.cutoff_lut\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_80_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_149_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08962_ channels.freq2\[9\] _01425_ _01290_ channels.freq1\[9\] _01426_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_110_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13668__A1 _04578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08893_ channels.accum\[0\]\[4\] _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__15715__I _07635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09713__I _01780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12891__A2 _04896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09514_ _01783_ _01826_ _01839_ _01905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_91_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12643__A2 _04537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09445_ _01788_ _01836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_140_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_140_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09376_ _01775_ _01776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_163_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14148__A2 _06016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_172_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12159__A1 _03317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08999__I _01460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10220_ _01509_ _02473_ _02480_ _02432_ _02481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_162_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15648__A2 _07579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10151_ channels.pw1\[8\] _01285_ _02412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10082_ _02348_ _02349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_50_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13910_ _05829_ _05910_ _05911_ _05912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_14890_ _06760_ _06869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16073__A2 _07924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10893__A1 _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13841_ _05811_ _05813_ _05843_ _05844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_57_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15820__A2 _07697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16560_ _08338_ _08340_ _00751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13772_ _05774_ _05775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12634__A2 _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10984_ _03201_ _03205_ _03209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_15511_ _07452_ _07453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_168_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12723_ _04477_ _04729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_84_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16491_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[2\] _08282_ _08252_ _08283_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15442_ net36 _07388_ _07389_ _07390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12654_ _04655_ _04657_ _04659_ _04660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_65_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12398__A1 _03398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11605_ _03675_ _03703_ _03708_ _00428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_38_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12585_ _04587_ _04589_ _04590_ _04591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_15373_ _07324_ _07325_ _07326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_37_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10948__A2 _01261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17112_ _00182_ clknet_leaf_116_clk channels.sus_rel1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_136_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11536_ _03639_ _03658_ _03661_ _00406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14324_ _06320_ _06321_ _06322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_68_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17043_ _00113_ clknet_leaf_225_clk channels.lfsr\[1\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14255_ _05560_ _06254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11467_ _03617_ _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_151_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13206_ _04277_ _04817_ _05212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10418_ _02677_ _02678_ _02679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_14186_ _01821_ _06186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_11398_ _03566_ _01487_ _03576_ _00353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13137_ _04389_ _04817_ _05143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_103_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10349_ _02597_ _02605_ _02610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12224__I _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13068_ _04926_ _05074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14311__A2 _06229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12322__A1 _04319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12019_ _04025_ _04076_ _04083_ _00467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_174_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_144_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16827_ tt_um_rejunity_sn76489.noise\[0\].gen.restart_noise _04158_ _00924_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16794__C _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16758_ _08453_ _00868_ _00874_ _00808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08829__B2 channels.freq1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_122_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15709_ _07630_ _07631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_75_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_88_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16689_ _08333_ _08429_ _08430_ _08431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_159_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09230_ channels.lfsr\[3\]\[11\] _01667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_173_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15575__A1 filters.sample_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12389__A1 _03381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09161_ _01601_ _01602_ _01594_ _01603_ _01605_ _01607_ _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_56_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15327__A1 filters.low\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09092_ channels.accum\[0\]\[19\] _01461_ _01546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_160_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09006__A1 channels.freq2\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14614__I _06186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09006__B2 channels.freq1\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_168_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09557__A2 _01899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12156__A4 filters.high\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09994_ channels.ctrl_reg3\[6\] _02283_ _02284_ _02287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_164_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08945_ _01400_ _01401_ _01410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_181_3743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11973__I _04011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08876_ _01345_ _01346_ _01347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09443__I _01833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09190__B1 _01632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_168_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16276__I _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09428_ filters.mode_vol\[7\] _01803_ _01809_ _01820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09359_ _01760_ _01761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_164_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12309__I _04314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13041__A2 _04991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11052__A1 filters.high\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12370_ _04375_ _04376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_63_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11321_ _01805_ _03492_ _03519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xclkbuf_5_16__f_clk clknet_3_4_0_clk clknet_5_16__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14040_ _06036_ _06040_ _06041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_105_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11252_ _03453_ _03392_ _03393_ _03462_ _00321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_24_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10203_ _01249_ _02427_ channels.pw3\[1\] _02464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_28_1193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11183_ _03397_ _03398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_10134_ _02360_ _02394_ _02395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_24_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15991_ spi_dac_i.spi_dat_buff_1\[0\] _07867_ _07870_ spi_dac_i.spi_dat_buff_1\[1\]
+ _07871_ _07872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_140_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_89_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17730_ _00800_ clknet_leaf_64_clk tt_um_rejunity_sn76489.control_tone_freq\[1\]\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_89_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10065_ filters.cutoff_lut\[11\] _02332_ _02335_ _02338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14942_ _05534_ _06915_ _06916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09353__I net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17661_ _00731_ clknet_leaf_81_clk tt_um_rejunity_sn76489.noise\[0\].gen.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14873_ filters.low\[26\] _06472_ _03473_ _06853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_16612_ _08374_ _08380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_173_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13824_ _05725_ _05736_ _05826_ _05827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_17592_ _00662_ clknet_leaf_38_clk spi_dac_i.spi_dat_buff_0\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12607__A2 _04566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_67_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16543_ _08324_ _08325_ _08313_ _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_58_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10967_ filters.filter_step\[1\] _03192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_13755_ _05752_ _05755_ _05758_ _05759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_168_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12706_ _04711_ _04712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_169_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16474_ _08241_ _08267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_100_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10898_ _02366_ _02831_ _03145_ _00284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13686_ filters.high\[22\] filters.band\[22\] _05179_ _05690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_182_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15425_ _07363_ _06862_ _07374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_38_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12637_ _04642_ _04643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_80_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12568_ _04563_ _04572_ _04573_ _04574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_15356_ filters.high\[19\] _07310_ _07223_ _07311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_170_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10397__A3 _02569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12791__A1 _04792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_152_Right_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_135_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11519_ _03641_ _03649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14307_ _06257_ _06272_ _06270_ _06305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_180_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12499_ _04406_ _04505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15287_ _03439_ _07231_ _07247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17026_ _00003_ clknet_leaf_240_clk filters.res_lut\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14238_ filters.band\[26\] _04596_ _06237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16809__A1 _08453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10149__A3 channels.pw2\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12543__A1 _04356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14169_ _05967_ _06062_ _06169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_146_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08730_ _01213_ _01214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_1_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08661_ _01144_ _01145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_1_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14048__A1 _04377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08592_ channels.lfsr\[3\]\[0\] _01107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_120_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13271__A2 _05188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11282__A1 _02316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10085__A2 _01905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09213_ channels.lfsr\[2\]\[10\] _01652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09144_ channels.lfsr\[2\]\[0\] _01593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11034__A1 filters.high\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11968__I _04006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08986__B1 _01448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09075_ channels.accum\[0\]\[17\] _01334_ _01530_ _01255_ _01531_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_86_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_135_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15720__A1 _05647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12534__A1 _04537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12799__I _04804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09977_ _02274_ _02276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08928_ _01337_ _01393_ _01394_ _01395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_157_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08859_ _01324_ _01330_ _01331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11870_ _03768_ _03957_ _03958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_19_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10821_ _03025_ _03042_ _03075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11273__A1 _03243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10752_ _02986_ _03007_ _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_13540_ _05544_ _05545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_149_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_9_Left_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13471_ _05313_ _05319_ _05476_ _05477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10683_ _02939_ _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_152_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12422_ _04364_ _04413_ _04427_ _04428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_15210_ _06918_ _07173_ _00568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_180_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16190_ _08061_ _08063_ _08042_ _08064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12773__A1 filters.cutoff_lut\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12353_ _04356_ _04358_ _04359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_15141_ _01760_ channels.sample2\[7\] _07107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09348__I _01750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11304_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[0\] _03506_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_65_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15072_ _07015_ _07038_ _07039_ _07040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12284_ _04273_ _04290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_22_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14023_ _05918_ _05934_ _06023_ _06024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_31_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11235_ _03445_ _03447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_121_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11166_ _03381_ _03382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_140_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_179_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10117_ _02377_ _02378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_93_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15974_ _07850_ _07852_ _07854_ _07855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11097_ _03316_ _03317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_141_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17713_ _00783_ clknet_leaf_74_clk tt_um_rejunity_sn76489.tone\[0\].gen.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10048_ _02324_ _02320_ _02325_ _00254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14925_ _06898_ _06900_ _00556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_117_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17644_ _00714_ clknet_leaf_206_clk channels.ch3_env\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_14856_ filters.band\[24\] _03474_ _06838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13807_ _05792_ _05809_ _05810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_82_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17575_ _00645_ clknet_leaf_38_clk spi_dac_i.counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_82_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14787_ filters.band\[17\] _04160_ _06775_ _06776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11999_ channels.env_counter\[2\]\[13\] _04012_ _04069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16526_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[8\] _08263_ _08311_ _08312_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_42_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13738_ _05662_ _05741_ _05742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_85_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16457_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[5\] _08251_ _07700_ _08254_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13669_ _05587_ _05589_ _05672_ _05673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_155_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11016__A1 _01069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15408_ _07345_ _07353_ _07358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_16388_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[3\] _08198_ _08203_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_29__f_clk_I clknet_3_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15339_ filters.low\[17\] _07295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_123_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14505__A2 _06501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09900_ channels.atk_dec2\[5\] _02220_ _02217_ _02222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_17009_ _00088_ clknet_leaf_225_clk channels.lfsr\[2\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09831_ channels.freq2\[13\] _02171_ _02167_ _02173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_130_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09762_ _02124_ _02125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09145__B1 _01592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08713_ _01191_ _01196_ _01197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_179_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09693_ channels.freq1\[8\] _02075_ _02036_ _02076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09696__A1 channels.freq1\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer11 _05431_ net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15723__I _07639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08644_ channels.env_vol\[3\]\[3\] _01133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer22 _06304_ net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer33 _05475_ net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15769__A1 _03468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_159_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08575_ _01091_ _00011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_107_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_176_3642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_176_3653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14992__A2 channels.sample1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09127_ channels.lfsr\[3\]\[17\] _01576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_115_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16497__A2 _08282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09058_ channels.accum\[0\]\[15\] _01461_ _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12507__A1 _04512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16503__B _08292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11020_ _03244_ _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_38_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14958__B _06921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12971_ _04808_ _04809_ _04977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_99_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09231__S0 _01305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14680__A1 filters.band\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14710_ _06703_ _06691_ _06704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_4
X_11922_ _04004_ _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_87_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15690_ _07615_ _07617_ _07618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14641_ _06619_ _06622_ _06635_ _06636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_157_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11853_ _03743_ _03939_ _03943_ _00441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_129_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14432__A1 _04802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17360_ _00430_ clknet_leaf_89_clk channels.pw2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10804_ _03038_ _03040_ _03058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_11784_ _03873_ _03874_ _03875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14572_ _04326_ _05891_ _06568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16311_ channels.env_counter\[3\]\[11\] _08153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_60_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13523_ _05293_ _05376_ _05529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10735_ _02953_ _02957_ _02991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_17291_ _00361_ clknet_leaf_189_clk channels.accum\[2\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16242_ spi_dac_i.spi_dat_buff_1\[11\] _07870_ _07700_ _08113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13454_ _05305_ _05320_ _05460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10666_ _02505_ _02923_ _02924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12405_ _04331_ _04338_ _04411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16173_ _08045_ _08023_ _08047_ _08048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13385_ _05382_ _05385_ _05390_ _05391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_97_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09611__A1 channels.pw2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10597_ _02850_ _02855_ _02856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__09611__B2 channels.freq2\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15124_ _07055_ _07059_ _07090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_11_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12336_ _04341_ _04342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_58_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12267_ _04272_ _04273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15055_ _07023_ _07024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_75_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14006_ _04742_ _05588_ _06007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11218_ filters.sample_filtered\[12\] _03430_ _03431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_43_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12198_ _04193_ _04202_ _04204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_177_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11149_ _03359_ _03230_ _03365_ _03366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_15957_ _07722_ _07838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_179_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09678__A1 filters.mode_vol\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14908_ _06718_ _06884_ _06885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__10288__A2 _02377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15888_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[0\] _07768_ _07770_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17627_ _00697_ clknet_leaf_208_clk channels.env_vol\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14839_ filters.low\[23\] _06822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__13226__A2 _05229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17558_ _00628_ clknet_leaf_244_clk filters.low\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16509_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[5\] _08289_ _08296_ _08297_
+ _08298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_119_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17489_ _00559_ clknet_leaf_13_clk filters.high\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_154_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_171_3550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_171_3561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09602__A1 filters.cutoff_lut\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10212__A2 _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09814_ _02160_ _02151_ _02161_ _00184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09118__B1 _01568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09745_ channels.ctrl_reg1\[2\] _02108_ _02113_ _02114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_158_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09676_ channels.sus_rel3\[7\] _01963_ _01964_ channels.sus_rel1\[7\] _02059_ _02060_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_119_1168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08627_ _01124_ _00030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_96_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08558_ _01074_ _01075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14965__A2 channels.sample3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08489_ filters.res_filt\[4\] _01005_ _01018_ _01019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__09841__A1 _02088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16706__A3 _03494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10520_ _02741_ _02780_ _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_174_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10451__A2 _02527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14717__A2 _06397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_99_Left_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10451_ _02508_ _02527_ _02712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_162_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13170_ _04703_ _04490_ _05176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10382_ _02642_ _02555_ _02643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12121_ _04142_ _00510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_130_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15142__A2 channels.sample1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_103_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13153__A1 _05158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12052_ _01063_ clk_ctr\[1\] _04102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12900__A1 _04895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11003_ _03207_ _03228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_53_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16860_ _03745_ _03775_ _00948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_53_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15811_ _06867_ _07698_ _07706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_102_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16791_ _07841_ _00899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09204__S0 _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_29_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15742_ _07332_ _07657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12954_ _04957_ _04958_ _04960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09361__I _01752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11905_ _03860_ _03861_ _03883_ _03988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_15673_ filters.sample_buff\[12\] _03450_ _07602_ _07603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_59_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12885_ _04886_ _04890_ _04891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14405__A1 _03361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_193_clk clknet_5_23__leaf_clk clknet_leaf_193_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_158_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17412_ _00482_ clknet_leaf_86_clk clk_ctr\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14624_ _06520_ _04601_ _06619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11836_ _03924_ _03925_ _03927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_114_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14956__A2 _06915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17343_ _00413_ clknet_leaf_102_clk channels.freq2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14555_ _06462_ _06463_ _06550_ _06551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09832__A1 _02155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11767_ _03857_ _03858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_138_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13506_ _04467_ _05512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_17274_ _00344_ clknet_leaf_186_clk channels.accum\[2\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10718_ _02974_ _02975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14708__A2 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14486_ _06354_ _06481_ _06482_ _06483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_11698_ channels.atk_dec1\[0\] channels.sus_rel1\[0\] _03784_ _03789_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_71_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12719__A1 _04458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16225_ _07683_ _08098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_70_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13437_ _05338_ _05355_ _05443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_36_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10649_ _02899_ _02906_ _02907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xrebuffer2 _05037_ net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__15381__A2 _07033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11131__I _03348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16156_ _08026_ _08028_ _08031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_141_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13368_ _05360_ _05364_ _05373_ _05374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_23_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15107_ _01760_ channels.sample2\[6\] _07074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12319_ _04324_ _04325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16087_ _07964_ _07936_ _07965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13299_ _05217_ _05224_ _05304_ _05305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_110_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15038_ _07001_ _07003_ _07006_ _07007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09899__A1 _02150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16989_ _00068_ clknet_leaf_164_clk channels.accum\[0\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_155_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09530_ channels.ch3_env\[1\] _01877_ _01920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09461_ filters.cutoff_lut\[6\] _01849_ _01851_ filters.cutoff_lut\[9\] _01852_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__11306__I _03507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09392_ _01790_ _01791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_3601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09823__A1 channels.freq2\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11630__A1 _03675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15372__A2 _07321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11933__A2 _03874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16321__A1 _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_35_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14635__A1 _05624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09728_ _01062_ _02100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_69_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09659_ channels.freq3\[6\] _01871_ _01999_ channels.ctrl_reg3\[6\] _02044_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_175_clk clknet_5_18__leaf_clk clknet_leaf_175_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_167_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12670_ _04560_ _04676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_38_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_207_clk_I clknet_5_20__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12949__A1 _04475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11621_ _03711_ _03719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_93_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09814__A1 _02160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14340_ _04326_ _05585_ _06338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11552_ _02154_ _03673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_80_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10503_ _02646_ _02647_ _02764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_150_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11483_ _03624_ _03625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14271_ _06259_ _06269_ _06270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_80_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16010_ _07775_ _07890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12177__A2 _04182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10434_ _02683_ _02693_ _02694_ _02695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13222_ _05227_ _05226_ _05228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_122_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10188__A1 channels.pw1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15358__I _07030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10365_ _02618_ _02625_ _02626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13153_ _05158_ _04510_ _05159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_55_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14262__I _06008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09356__I filters.filt_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12104_ channels.accum\[3\]\[0\] _04134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_72_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13084_ _05076_ _05088_ _05089_ _05090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10296_ _01307_ _02556_ _02557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_72_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12035_ _04051_ _04090_ _04093_ _00473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16912_ _00985_ _00851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11688__A1 _03534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08553__A1 channels.clk_div\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11783__S1 _01167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16843_ _00932_ _00933_ _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10360__A1 _01542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16774_ _03499_ _00886_ _00887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13986_ _05985_ _05986_ _05987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_88_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15725_ _03268_ _07643_ _07644_ _07645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_125_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10112__A1 channels.ctrl_reg2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12937_ _04863_ _04865_ _04943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xclkbuf_leaf_166_clk clknet_5_25__leaf_clk clknet_leaf_166_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_38_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15656_ filters.sample_buff\[10\] _07579_ _07587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_12868_ _04871_ _04872_ _04873_ _04874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_69_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14607_ _06400_ _06502_ _06603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_103_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11819_ _03906_ _03847_ _03909_ _03910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_133_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15042__B _04993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15587_ _07449_ _07523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12799_ _04804_ _04805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13341__I _05259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17326_ _00396_ clknet_leaf_87_clk channels.freq1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14538_ _06523_ _06533_ _06534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_138_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17257_ _00327_ clknet_leaf_71_clk tt_um_rejunity_sn76489.control_tone_freq\[0\]\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__16551__A1 _08314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14469_ _06460_ _06465_ _06466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16208_ _08064_ _08067_ _08081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13365__A1 _04641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17188_ _00258_ clknet_leaf_79_clk filters.cutoff_lut\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_11_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11376__B1 _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16139_ _08014_ _07961_ _07858_ _08015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15106__A2 channels.sample3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_149_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16854__A2 _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08961_ _01276_ _01425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_166_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13668__A2 _05671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_166_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_166_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11679__A1 channels.sus_rel2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11679__B2 channels.sus_rel1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08892_ _01322_ _01359_ _01361_ _00058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_127_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09513_ _01903_ _01904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_151_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_157_clk clknet_5_29__leaf_clk clknet_leaf_157_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_91_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09444_ channels.ctrl_reg2\[0\] _01830_ _01834_ channels.freq3\[8\] _01835_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_140_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_166_Right_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_74_Right_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_176_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09375_ net11 _01775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_136_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11603__A1 _03673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17250__CLK clknet_5_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_193_clk_I clknet_5_23__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_5_0_clk clknet_0_clk clknet_3_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_171_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_73_clk_I clknet_5_14__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_83_Right_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_101_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10150_ _02389_ _02405_ channels.pw3\[8\] _02411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14856__A1 filters.band\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_88_clk_I clknet_5_12__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10081_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[4\] tt_um_rejunity_sn76489.noise\[0\].gen.counter\[5\]
+ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[6\] _02347_ tt_um_rejunity_sn76489.control_noise\[0\]\[0\]
+ tt_um_rejunity_sn76489.control_noise\[0\]\[1\] _02348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_131_clk_I clknet_5_31__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12882__A3 _04803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13840_ _05825_ _05842_ _05843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_11_clk_I clknet_5_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10893__A2 _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_148_clk clknet_5_31__leaf_clk clknet_leaf_148_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13771_ _05687_ _05774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_58_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10983_ filters.low\[0\] _03188_ _03200_ _03207_ _03208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA_clkbuf_leaf_146_clk_I clknet_5_28__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_92_Right_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15510_ _03202_ _03204_ _03215_ _07452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_12722_ _04236_ _04728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16490_ _08281_ _08282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_57_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_133_Right_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15441_ _07373_ _07370_ _07376_ _07374_ _07389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA_clkbuf_leaf_26_clk_I clknet_5_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12653_ _04658_ _04639_ _04659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_182_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16781__A1 _02098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_65_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11604_ channels.pw3\[6\] _03704_ _03705_ _03708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12398__A2 _04403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13595__A1 _05591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15372_ _07315_ _07321_ _07325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_182_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12584_ _04560_ _04586_ _04559_ _04590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_182_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17111_ _00181_ clknet_leaf_114_clk channels.sus_rel1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_167_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14323_ _04858_ _05487_ _06321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11535_ channels.freq2\[0\] _03659_ _03660_ _03661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16533__A1 _08314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17042_ _00112_ clknet_leaf_226_clk channels.lfsr\[1\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14254_ _06194_ _06252_ _06253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_34_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11466_ channels.accum\[1\]\[17\] _01230_ _01530_ _01101_ _03617_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_21_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13205_ _05143_ _05209_ _05210_ _05211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10417_ _02655_ _02630_ _02641_ _02678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_14185_ _05975_ _06184_ _06185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11397_ channels.accum\[2\]\[13\] _03571_ _03576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09086__I _01321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16836__A2 _03731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13136_ _05139_ _05140_ _05141_ _05142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_10348_ _02548_ _02563_ _02608_ _02609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__10025__I _02104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13067_ _05066_ _05072_ _05073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10279_ _01470_ _02539_ _02540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_40_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08526__A1 _01043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12322__A2 _04327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12018_ channels.env_counter\[1\]\[3\] _04079_ _04083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_144_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16064__A3 _07942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16826_ _03490_ _00922_ _03519_ _00923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_136_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16757_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[6\] _00873_ _00871_ _00874_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_139_clk clknet_5_31__leaf_clk clknet_leaf_139_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13969_ _03299_ _03471_ _05970_ _05971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_122_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15708_ _07629_ _07630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_75_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16688_ _08425_ _08428_ _08430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_61_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15639_ _07486_ _07570_ _07571_ _07572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_100_Right_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_150_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15575__A2 _07504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09160_ _01606_ _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12389__A2 _04341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_173_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17309_ _00379_ clknet_leaf_158_clk channels.accum\[1\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_173_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09091_ _01449_ _01544_ _01545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13338__A1 _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_168_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_168_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16827__A2 _04158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12561__A2 _04566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09993_ _02238_ _02282_ _02286_ _00238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10572__A1 channels.sample3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08944_ _01257_ _01409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_122_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08517__A1 _01043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_181_3744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12313__A2 _04318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08875_ _01343_ _01346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_93_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_4_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input15_I bus_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09493__A2 _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09427_ _01818_ _01819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_176_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13577__A1 _05508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09358_ _01759_ _01760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_62_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_43_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09289_ channels.lfsr\[2\]\[22\] _01716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11320_ _03515_ _03508_ _03518_ _00333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_133_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11251_ _03454_ _03461_ _03462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_120_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_26_Left_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10202_ _01469_ _02460_ _02461_ _02462_ _02463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_31_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11182_ _03247_ _03379_ _03250_ _03396_ _03397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_101_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10133_ _02391_ _02392_ _02393_ _02394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_15990_ _02101_ _07871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_89_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10064_ _02314_ _02331_ _02337_ _00258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14941_ _04558_ _04690_ _06915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_89_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17660_ _00730_ clknet_leaf_82_clk tt_um_rejunity_sn76489.noise\[0\].gen.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14872_ _06706_ _06852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16611_ _01615_ _08376_ _08379_ _01617_ _00763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_13823_ _05728_ _05735_ _05826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17591_ _00661_ clknet_leaf_42_clk spi_dac_i.spi_dat_buff_1\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_35_Left_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_67_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16542_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[0\] _08263_ _08325_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13754_ _05537_ _05756_ _05757_ _05758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_15_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10966_ _03190_ _03191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_57_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12705_ filters.high\[12\] filters.band\[12\] _04710_ _04711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_16473_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[1\] _08266_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13685_ _04294_ _05260_ _05689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10897_ channels.sample2\[1\] _03143_ _03145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_100_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15424_ _07372_ _07373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__13568__A1 _04764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12636_ _04641_ _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_171_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12240__A1 _04233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15355_ _07029_ _07310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12567_ _04570_ _04571_ _04573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_26_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14306_ _05877_ _06300_ _06302_ _06303_ _06304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_11518_ _03515_ _03642_ _03648_ _00401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12791__A2 _04796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15286_ _05968_ _07245_ _07246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12498_ _04201_ _04504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_44_Left_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17025_ _00002_ clknet_leaf_240_clk filters.res_lut\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14237_ _06234_ _06235_ _06236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_151_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11449_ channels.accum\[1\]\[10\] _03607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_180_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14168_ _06164_ _06167_ _06168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_42_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13119_ _05123_ _05124_ _05125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_14099_ _06092_ _06098_ _06099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09544__I _01932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input7_I bus_cyc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08660_ _01143_ _01144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_1_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14048__A2 _05074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_53_Left_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16809_ _08453_ _00906_ _00911_ _00910_ _00822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_72_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08591_ _01106_ _00012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_17789_ _00859_ clknet_leaf_49_clk tt_um_rejunity_sn76489.control_noise\[0\]\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_3_4_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_5_22__f_clk clknet_3_5_0_clk clknet_5_22__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_163_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16745__A1 _01800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15548__A2 _07478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13559__A1 _05563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09212_ _01646_ _01634_ _01650_ _01651_ _00088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_63_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09143_ _01591_ _01592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_173_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_62_Left_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09719__I _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09074_ _01323_ _01529_ _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_112_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_20_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15720__A2 _07640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09976_ _02274_ _02275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_110_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14287__A2 _06285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08927_ _01385_ _01386_ _01392_ _01394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XPHY_EDGE_ROW_71_Left_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08858_ _01327_ _01329_ _01330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_58_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08789_ _01261_ _01262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15787__A2 _07682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13798__A1 _05512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10820_ _03058_ _03073_ _03074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_39_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10751_ _02987_ _03006_ _03007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_67_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15539__A2 _07478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13470_ _05307_ _05312_ _05476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_62_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10682_ _02923_ _02939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_168_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_80_Left_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_125_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12421_ _04415_ _04419_ _04426_ _04427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_36_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_164_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08977__A1 channels.freq3\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15140_ _01770_ channels.sample3\[7\] _07106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12352_ _04357_ _04249_ _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_65_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13970__A1 _05968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11303_ _02299_ _03498_ _03505_ _00329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__16750__I _00867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12055__I _04103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15071_ _07017_ _07021_ _07039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_12283_ _04206_ _04288_ _04289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14022_ _05920_ _05933_ _06023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13722__A1 _05631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11234_ _03436_ _03438_ _03445_ _03446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_120_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_8_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11165_ _03247_ _03379_ _03250_ _03380_ _03381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XANTENNA__09364__I net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10116_ _02360_ _02376_ _02377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_15973_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[1\] _07853_ _07854_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11096_ _03315_ _03316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_141_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10047_ channels.sus_rel3\[5\] _02321_ _02322_ _02325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_17712_ _00782_ clknet_leaf_218_clk channels.lfsr\[0\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14924_ filters.band\[30\] _06869_ _06899_ _06900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_136_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14855_ filters.low\[24\] _06837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_17643_ _00713_ clknet_leaf_206_clk channels.ch3_env\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_37_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13806_ _05799_ _05808_ _05809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_17574_ _00644_ clknet_leaf_6_clk filters.filter_step\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XTAP_TAPCELL_ROW_82_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14786_ _03721_ _06775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_11998_ _04044_ _04067_ _04068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_82_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16525_ _08238_ _08305_ _08309_ _08311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_9_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13737_ _05678_ _05681_ _05740_ _05741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_46_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10949_ _03174_ _03122_ _03176_ _00304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_27_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_70_clk clknet_5_14__leaf_clk clknet_leaf_70_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_2_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16456_ _08251_ _08253_ _00734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13668_ _04578_ _05671_ _05590_ _05672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_42_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_155_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15407_ _07312_ _07354_ _07357_ _00581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_26_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12619_ _04623_ _04624_ _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_16387_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[2\] _08201_ _08202_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_182_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13599_ net62 _05492_ _05603_ _05604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_14_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12764__A2 _04766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15338_ _07280_ _07284_ _07294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_117_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10775__A1 _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15269_ _07206_ _07228_ _07229_ _07230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_111_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17008_ _00087_ clknet_leaf_222_clk channels.lfsr\[2\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09393__A1 _01781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09830_ _02150_ _02170_ _02172_ _00189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_21_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_130_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09761_ _02123_ _01901_ _02124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08712_ _01174_ _01192_ _01195_ _01196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09692_ _02073_ _02075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xrebuffer12 _05060_ net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_179_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xrebuffer23 _04988_ net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08643_ _01132_ _00038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer34 _03286_ net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15769__A2 _07670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08574_ _01084_ _01086_ _01090_ channels.ring_outs\[2\] _01091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09448__A2 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_176_3643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_176_3654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_61_clk clknet_5_9__leaf_clk clknet_leaf_61_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_9_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_76_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_137_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08959__A1 _01414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09126_ channels.lfsr\[2\]\[17\] _01575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09057_ _01449_ _01514_ _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11928__B _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09959_ channels.freq3\[15\] _02258_ _02262_ _02263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12970_ _04448_ _04461_ _04976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__15209__A1 filters.high\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09231__S1 _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11921_ _04001_ _04003_ _04004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__13434__I _04562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14640_ _06627_ _06628_ _06634_ _06635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_11852_ channels.env_vol\[0\]\[0\] _03942_ _03943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10803_ _03055_ _03056_ _03057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14571_ _06426_ _06427_ _06566_ _06567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_11783_ channels.env_counter\[0\]\[1\] channels.env_counter\[1\]\[1\] channels.env_counter\[2\]\[1\]
+ channels.env_counter\[3\]\[1\] _03831_ _01167_ _03874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
Xclkbuf_leaf_52_clk clknet_5_10__leaf_clk clknet_leaf_52_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_138_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16310_ _08152_ _00689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13522_ _05295_ _05528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_60_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10734_ _02988_ _02989_ _02990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17290_ _00360_ clknet_leaf_158_clk channels.accum\[2\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16241_ spi_dac_i.spi_dat_buff_1\[10\] _07722_ _08111_ _08107_ _08112_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_125_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13453_ _05457_ _05357_ _05458_ _05459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_10665_ _02768_ _02920_ _02922_ _02774_ _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_82_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12404_ _04409_ _04410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_16172_ _08046_ _08047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_24_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13384_ _05388_ _05389_ _05390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10596_ _02851_ _02854_ _02855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_97_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15123_ _03343_ _07064_ _07088_ _07089_ _00565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_11_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12335_ _03238_ _03182_ _04188_ _03373_ _04341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_133_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_146_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15054_ filters.low\[5\] _07022_ _07023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_118_Left_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12266_ _03362_ _04271_ _04272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_120_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14005_ _04529_ _06005_ _06006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_75_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11217_ _03426_ _03429_ _03430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11801__S0 _03886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12197_ _04193_ _04202_ _04203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_37_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11148_ _03360_ _03220_ _03364_ _03344_ _03365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_37_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15956_ _07598_ _07837_ _00650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11079_ _03246_ _03283_ _03249_ _03299_ _03300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_37_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13474__A3 _04804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14907_ _06882_ _03475_ _06883_ _06884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_15887_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[1\] _07766_ _07769_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_17626_ _00696_ clknet_leaf_209_clk channels.env_vol\[1\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_127_Left_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_114_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14838_ _06819_ _06821_ _00548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_148_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14769_ _06748_ _06758_ _06759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_17557_ _00627_ clknet_leaf_27_clk filters.low\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16508_ _08291_ _08295_ _08292_ _08297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17488_ _00558_ clknet_leaf_13_clk filters.high\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_160_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_154_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_154_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16439_ _08235_ _08236_ _08240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_143_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_171_3551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_171_3562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12737__A2 _04742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13934__A1 _05803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_132_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_111_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09813_ channels.sus_rel1\[7\] _02152_ _02158_ _02161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10920__A1 channels.sample2\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14111__A1 _03413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09744_ _02093_ _02113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_94_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09669__A2 net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09675_ _01908_ _02055_ _02057_ _02058_ _02059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_69_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_179_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13254__I _05259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08626_ channels.lfsr\[3\]\[17\] _01124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14414__A2 _06370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08557_ _01073_ _01074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13622__B1 _05626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_34_clk clknet_5_2__leaf_clk clknet_leaf_34_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_37_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08488_ _01017_ _01005_ _01018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09841__A2 _01862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14178__A1 _03329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10450_ _02505_ _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__10739__A1 _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16514__B _08301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09109_ channels.accum\[0\]\[21\] _01560_ _01561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10381_ _02641_ _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10203__A3 channels.pw3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15678__A1 _07598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12120_ channels.accum\[3\]\[8\] _04142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12051_ _02353_ _04101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_92_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11002_ filters.lp _03226_ _03227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12900__A2 _04900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14102__A1 _06024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15810_ _07704_ _07705_ _00636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16790_ _00892_ _00896_ _00898_ _00889_ _00816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_70_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09204__S1 _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15741_ _07639_ _07656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12953_ _04957_ _04958_ _04959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_29_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11904_ _03930_ _03904_ _03908_ _03986_ _03987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_87_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15672_ _07601_ _07602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12884_ _04887_ _04888_ _04889_ _04890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__13208__A3 _05106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17411_ _00481_ clknet_leaf_86_clk clk_ctr\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14623_ _04222_ _06383_ _06618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11835_ _03924_ _03925_ _03926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_leaf_25_clk clknet_5_6__leaf_clk clknet_leaf_25_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_17342_ _00412_ clknet_leaf_100_clk channels.freq2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14554_ _06359_ _06093_ _06464_ _06550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_99_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11766_ _03815_ _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_55_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13505_ _05509_ _04758_ _04946_ _05510_ _05511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__14169__A1 _05967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17273_ _00343_ clknet_leaf_179_clk channels.accum\[2\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10717_ _01088_ _02974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_125_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14485_ _06355_ _06357_ _06482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_11697_ _01290_ _03788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_125_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09089__I _01542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16224_ spi_dac_i.spi_dat_buff_1\[8\] _07834_ _08093_ _08095_ _08096_ _08097_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_125_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12719__A2 _04459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13436_ _05369_ _05371_ _05441_ _05442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_64_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10648_ _02904_ _02905_ _02906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09045__B1 _01503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrebuffer3 net42 net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_77_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16155_ _07743_ _08029_ _08030_ _00656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_77_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13367_ _05365_ _05372_ _05373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_106_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14723__I _06703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10579_ _02687_ _02777_ _02817_ _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_106_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15669__A1 filters.sample_buff\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15106_ _01769_ channels.sample3\[6\] _07073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12318_ _04323_ _04324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16086_ _07931_ _07964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13298_ _05211_ _05216_ _05304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_110_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14341__A1 _04378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15037_ _06997_ _07000_ _07006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_12249_ _04254_ _04255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_120_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10902__A1 channels.sample2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16094__A1 _07929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08571__A2 _01083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16988_ _00067_ clknet_leaf_151_clk channels.accum\[0\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_147_Right_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15939_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[1\] _07821_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_78_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09520__A1 _01823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09460_ _01000_ _01850_ _01851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_64_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17609_ _00679_ clknet_leaf_131_clk channels.env_counter\[3\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_171_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09391_ _01783_ _01785_ _01789_ _01790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_19_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_173_3602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_15_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09587__A1 channels.pw1\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_13__f_clk_I clknet_3_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11394__A1 _03566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10197__A2 _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16321__A2 _03936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_35_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_114_Right_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14635__A2 _05281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09727_ _02098_ _02091_ _02099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09511__B2 channels.atk_dec1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10401__I _02561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09658_ channels.pw2\[6\] _01996_ _01997_ channels.freq2\[14\] _02043_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_85_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08609_ _01115_ _00021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_38_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09589_ channels.sample3\[7\] _01977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_139_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11620_ _03666_ _03712_ _03718_ _00433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_37_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12949__A2 _04482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11551_ _03668_ _03669_ _03672_ _00410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_53_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10502_ _02744_ _02762_ _02763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_52_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14270_ _06267_ _06268_ _06269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11482_ _02289_ _01954_ _03624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_18_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13221_ _05159_ _05162_ _05227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_94_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10433_ _02669_ _02670_ _02666_ _02694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_13152_ _04366_ _05158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_66_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10364_ _02504_ _02624_ _02625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_55_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12103_ _04133_ _00501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14323__A1 _04858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13083_ _05080_ _05081_ _05089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_72_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10295_ channels.ch3_env\[1\] _02556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_72_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12034_ channels.env_counter\[1\]\[9\] _04091_ _04093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16911_ channels.exp_counter\[3\]\[4\] _00985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12885__A1 _04886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08553__A2 _01069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16842_ tt_um_rejunity_sn76489.clk_counter\[2\] _00931_ _01753_ _00933_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_1308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15823__A1 _03735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09189__S0 _01141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16773_ _00884_ _00886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13985_ _05937_ _05957_ _05986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_5_3__f_clk clknet_3_0_0_clk clknet_5_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12936_ _04863_ _04865_ _04942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_15724_ _07332_ _07644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10112__A2 channels.ring_outs\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15655_ filters.sample_buff\[11\] _07448_ _07586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12867_ _04814_ _04870_ _04873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15051__A2 channels.sample1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11818_ channels.env_counter\[0\]\[12\] channels.env_counter\[1\]\[12\] channels.env_counter\[2\]\[12\]
+ channels.env_counter\[3\]\[12\] _01150_ _01166_ _03909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_14606_ _06599_ _06601_ _06602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_15586_ _07511_ _07522_ _07435_ _00595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13062__A1 _03398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12798_ _04803_ _04804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_173_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17325_ _00395_ clknet_leaf_99_clk channels.freq1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14537_ _06526_ _06532_ _06533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11749_ _03837_ _03839_ _03840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_138_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17256_ _00326_ clknet_leaf_73_clk tt_um_rejunity_sn76489.control_tone_freq\[0\]\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14468_ _06461_ _06464_ _06465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_141_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09569__A1 channels.atk_dec2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16207_ _07882_ _07887_ _08065_ _08080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09569__B2 channels.pw3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13419_ _05379_ _05403_ _05425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_180_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17187_ _00257_ clknet_leaf_78_clk filters.cutoff_lut\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_141_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14399_ _05853_ _06397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_84_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11376__B2 _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16138_ _07773_ _08014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13069__I _05074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13117__A2 _04315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16069_ _07926_ _07947_ _07948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08960_ channels.freq3\[9\] _01077_ _01424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_149_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_5_clk clknet_5_4__leaf_clk clknet_leaf_5_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_110_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_166_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_166_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08891_ channels.accum\[0\]\[3\] _01360_ _01361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16067__A1 _07880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09741__A1 channels.ctrl_reg1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_127_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14829__S _06073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09512_ _01783_ _01824_ _01785_ _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_91_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09443_ _01833_ _01834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_148_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_140_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_164_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09374_ _01767_ _01743_ _01774_ _00127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_19_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16542__A2 _08263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11367__B2 _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14305__A1 _06275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09980__A1 _02245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10080_ tt_um_rejunity_sn76489.chan\[2\].attenuation.in _02347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_50_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09192__I _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14608__A2 _06501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13770_ _04630_ _05766_ _05773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10982_ _03206_ _03207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09920__I _02226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12721_ _04723_ _04726_ _04727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_97_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15440_ _07366_ _07387_ _07388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_48_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12652_ _04636_ _04658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_167_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13044__A1 _04928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11603_ _03673_ _03703_ _03707_ _00427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_65_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12058__I _04106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15371_ _07313_ _07314_ _07324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12583_ _04583_ _04584_ _04588_ _04589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_0_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17110_ _00180_ clknet_leaf_114_clk channels.sus_rel1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14322_ _05469_ _06027_ _06320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11534_ _03651_ _03660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08471__A1 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17041_ _00111_ clknet_leaf_225_clk channels.lfsr\[1\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14253_ _06230_ _06251_ _06252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_20_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11465_ _03614_ _03615_ _01524_ _03616_ _00380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11358__A1 _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13204_ _04320_ _04368_ _04882_ _05145_ _05210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__09367__I filters.filt_3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10416_ _02655_ _02676_ _02600_ _02677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_21_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14184_ _06180_ _06183_ _06184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_11396_ _03575_ _03569_ _01475_ _03570_ _00352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_150_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10030__A1 channels.sus_rel3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09971__A1 _02098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13135_ _05105_ _05108_ _05141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_103_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10347_ _02502_ _02607_ _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13066_ _05071_ _05067_ _05072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_40_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10278_ _02378_ _02539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_104_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12017_ _04021_ _04076_ _04082_ _00466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09723__A1 channels.pw1\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_144_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11530__A1 _02328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16825_ _03496_ _00922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_161_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16756_ _00867_ _00873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_105_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13968_ _05969_ _03471_ _05970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_49_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_122_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15707_ _07443_ _03214_ _07628_ _07629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_12919_ _04175_ _04924_ _04925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_85_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_100_Left_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16687_ _08425_ _08428_ _08429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13899_ _05813_ _05843_ _05901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15638_ _07562_ _07557_ _07569_ _07571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_131_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_174_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15569_ _07499_ _07496_ _07506_ _07507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_145_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17308_ _00378_ clknet_leaf_154_clk channels.accum\[1\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09090_ _01537_ _01543_ _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_160_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15500__C _06917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13338__A2 _04739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17239_ _00309_ clknet_leaf_91_clk filters.sample_filtered\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11349__A1 _03535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_168_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_3_0_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16288__A1 _02354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08765__A2 _01090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12561__A3 _04504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09992_ channels.ctrl_reg3\[5\] _02283_ _02284_ _02286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_161_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08943_ channels.accum\[0\]\[8\] _01408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_206_clk_I clknet_5_22__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12849__A1 _03364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_181_3734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09714__A1 _02088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08517__A2 _01008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_181_3745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08874_ _01338_ _01332_ _01345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_1295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_4_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15742__I _07332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09740__I _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13262__I _05092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09426_ _01817_ _01818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_177_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14774__A1 filters.band\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09357_ _01758_ _01759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_164_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09288_ _01711_ _01591_ _01715_ _01699_ _00100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_43_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16515__A2 _08289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_43_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13329__A2 _05254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11250_ _03452_ _03460_ _03461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_120_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16279__A1 _08136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10012__A1 channels.atk_dec3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10201_ channels.pw1\[0\] _02435_ _02462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09953__A1 _02234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11181_ filters.band\[10\] _03396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_113_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10132_ channels.pw1\[11\] _01251_ _02393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_98_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09705__A1 _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17056__D _00126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10063_ filters.cutoff_lut\[10\] _02332_ _02335_ _02337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_89_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14940_ _06911_ _06912_ _06913_ _06914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_89_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11512__A1 _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14871_ _05546_ _06851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16610_ _01608_ _08376_ _08379_ _01612_ _00762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_13822_ _05816_ _05824_ _05825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_173_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17590_ _00660_ clknet_leaf_42_clk spi_dac_i.spi_dat_buff_1\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10079__A1 _02328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16541_ _08257_ _08323_ _08324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13753_ _05644_ _05645_ _05649_ _05757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_35_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10965_ _03189_ _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_85_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12704_ _03184_ _04710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_97_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16472_ _08135_ _08265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13684_ _04176_ _05687_ _05688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10896_ _02366_ _02783_ _03144_ _00283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_100_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15423_ filters.low\[25\] _07372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12635_ _04207_ _04641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13568__A2 _05570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15354_ _07305_ _07308_ _07309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_142_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12566_ _04570_ _04571_ _04572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_124_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12240__A2 _04245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11517_ channels.pw1\[3\] _03643_ _03644_ _03648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14305_ _06275_ _06277_ _06303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_80_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15285_ filters.low\[14\] _07244_ _07245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_135_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12497_ _04292_ _04288_ _04503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09097__I _01549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14236_ _06125_ _06133_ _06235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17024_ _00001_ clknet_leaf_240_clk filters.res_lut\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11448_ _03600_ _01433_ _03606_ _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09539__A4 _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09944__A1 channels.freq3\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08747__A2 _01105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14167_ _05977_ _06165_ _06166_ _06167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_104_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11379_ channels.accum\[2\]\[6\] _03565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_21_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13118_ _03332_ net60 _04450_ _05124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_14098_ _06095_ _06097_ _06098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13049_ _04641_ _05049_ _05055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12251__I _04218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11503__A1 channels.freq1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_179_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17240__CLK clknet_5_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_192_clk_I clknet_5_23__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16808_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[2\] _00907_ _00911_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08590_ _01086_ _01101_ _01105_ channels.ring_outs\[1\] _01106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_17788_ _00858_ clknet_leaf_56_clk tt_um_rejunity_sn76489.control_noise\[0\]\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_4_0_clk clknet_0_clk clknet_3_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_89_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_72_clk_I clknet_5_14__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16739_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[6\] _00861_ _08459_ _00862_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_159_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09211_ _01626_ _01651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16958__CLK clknet_5_16__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10490__A1 _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14756__A1 _05544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_87_clk_I clknet_5_12__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09142_ _01590_ _01591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_84_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_130_clk_I clknet_5_30__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09073_ _01526_ _01528_ _01529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_114_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_1254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_114_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_145_clk_I clknet_5_30__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09975_ _02208_ _01881_ _02274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_clkbuf_leaf_25_clk_I clknet_5_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08926_ _01385_ _01386_ _01392_ _01393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_58_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08857_ channels.accum\[0\]\[1\] channels.accum\[1\]\[1\] channels.accum\[2\]\[1\]
+ channels.accum\[3\]\[1\] _01307_ _01328_ _01329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_93_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15236__A2 _07168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_220_clk clknet_5_21__leaf_clk clknet_leaf_220_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08788_ _01256_ _01261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11505__I _01740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10750_ _02990_ _03005_ _03006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_39_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09409_ filters.lp _01803_ _01796_ _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10681_ _02917_ _02918_ _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_62_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12420_ _04421_ _04425_ _04426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_47_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_153_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08814__I _01286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12351_ _04252_ _04264_ _04283_ _04357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__12336__I _04341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11302_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[3\] _03500_ _03503_ _03505_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_121_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15172__A1 _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15070_ _07017_ _07021_ _07038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_121_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12282_ _04287_ _04288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_105_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14021_ _06002_ _06021_ _06022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09926__A1 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11233_ filters.sample_filtered\[13\] _03444_ _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13722__A2 _05632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10536__A2 _02754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11164_ filters.band\[9\] _03380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_8_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10115_ _02373_ _02374_ _02375_ _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_140_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15972_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[3\] _07790_ _07853_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_11095_ _03311_ _03312_ _03313_ _03314_ _03315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_41_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17711_ _00781_ clknet_leaf_231_clk channels.lfsr\[0\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_141_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10046_ _02154_ _02324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_117_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14923_ _06762_ _06899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_211_clk clknet_5_20__leaf_clk clknet_leaf_211_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_17642_ _00712_ clknet_leaf_206_clk channels.ch3_env\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_76_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14854_ _06701_ _06836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09380__I _01003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13805_ _05803_ _05807_ _05808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_86_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17573_ _00643_ clknet_5_5__leaf_clk filters.filter_step\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_11997_ _03920_ _04066_ _04067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_82_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14785_ _06771_ _06773_ _06774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_82_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16524_ _08280_ _08305_ _08309_ _08310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_86_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13736_ _05703_ _05705_ _05739_ _05740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_10948_ channels.sample1\[9\] _01261_ _03176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_27_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16455_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[4\] _08249_ _08252_ _08253_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13667_ _05585_ _05671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10879_ _03128_ _02890_ _03129_ _03130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_73_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15406_ filters.high\[23\] _07310_ _07356_ _07357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_38_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12618_ _04604_ _04605_ _04595_ _04624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_16386_ _08191_ _08201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13598_ _05477_ _05491_ _05603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13410__A1 _05405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12549_ _04551_ _04553_ _04555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_15337_ _07291_ _07292_ _07293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_108_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11972__A1 _04044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_152_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_1 _01588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15268_ _07210_ _07215_ _07229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_123_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09917__A1 channels.sus_rel2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17007_ _00086_ clknet_leaf_222_clk channels.lfsr\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14219_ _06129_ _06130_ _06218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_1_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15199_ filters.low\[10\] _05532_ _07162_ _07163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_67_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_130_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09760_ _01780_ _02123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08711_ _01179_ _01193_ _01194_ _01173_ _01195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_09691_ _02073_ _02074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_174_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_202_clk clknet_5_21__leaf_clk clknet_leaf_202_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08642_ channels.env_vol\[3\]\[2\] _01132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer13 net53 net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13229__A1 _04324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer24 net54 net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_178_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer35 net63 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_90_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08573_ _01089_ _01090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11335__S0 _01146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_176_3644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_176_3655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13540__I _05544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_137_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09125_ channels.lfsr\[1\]\[17\] _01574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10215__A1 _01541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10215__B2 _01533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08959__A2 _01415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16851__I _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11963__A1 _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15154__A1 _06913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09056_ _01512_ _01513_ _01514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11715__A1 channels.sus_rel3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11715__B2 channels.sus_rel2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09384__A2 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09958_ _02254_ _02262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_95_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08909_ _01375_ _01376_ _01377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09889_ channels.atk_dec2\[2\] _02211_ _02206_ _02214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15209__A2 _06934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11920_ _03534_ _04002_ _01585_ _04003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08895__A1 _01354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_1191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11851_ _03941_ _03942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_169_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_1164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_170_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10802_ _03015_ _03017_ _03051_ _03056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14570_ _04446_ _05449_ _06428_ _06566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11782_ _03871_ _03872_ _03873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13521_ _05435_ _05439_ _05526_ _05527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_0_32_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10733_ _02959_ _02967_ _02989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16240_ _08083_ _08104_ _08103_ _08111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13452_ _05303_ _05332_ _05458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10664_ _01085_ _02770_ _02921_ _02922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_12403_ _04383_ _04394_ _04408_ _04409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__10206__A1 _01481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16171_ _08017_ _08021_ _08046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13383_ _05382_ _05385_ _05389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_106_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10595_ _02852_ _02853_ _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_180_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_97_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12334_ _04291_ _04266_ _04340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15122_ _06186_ _07089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15053_ _07015_ _07017_ _07021_ _07022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_12265_ _03238_ _03203_ _04188_ _03359_ _04271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_121_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_128_Right_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_107_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09375__I net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14004_ _05943_ _06005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_75_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11216_ filters.high\[12\] _03428_ _03429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_112_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12196_ _03288_ _04197_ _04201_ _04202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_75_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11801__S1 _01170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16710__B _08318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11147_ _03363_ _03364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_128_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15955_ spi_dac_i.spi_dat_buff_1\[0\] _07728_ _07833_ _07836_ _07837_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_11078_ filters.band\[4\] _03299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_10029_ _02293_ _02312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14906_ _06456_ _03475_ _06883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08886__A1 _01354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15886_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[2\] _07765_ _07768_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_17625_ _00695_ clknet_leaf_209_clk channels.env_vol\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14959__A1 _06909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14837_ filters.band\[22\] _06820_ _06811_ _06821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17556_ _00626_ clknet_leaf_246_clk filters.low\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14768_ _06753_ _06757_ _06758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_16507_ _08291_ _08295_ _08296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10445__A1 _01162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13719_ _03398_ _04403_ _04805_ _05723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_73_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17487_ _00557_ clknet_leaf_23_clk filters.band\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14699_ _06602_ _06607_ _06693_ _06694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_154_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16438_ _08136_ _08239_ _00730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_26_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_171_3552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_171_3563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13934__A2 _05807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16369_ channels.ch3_env\[6\] _08185_ _08188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08810__A1 channels.ctrl_reg2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12704__I _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13698__A1 _05686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11173__A2 _03366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16636__A1 _01577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08574__B1 _01090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09812_ _01818_ _02160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_94_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10920__A2 _03156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09743_ _01766_ _02112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14111__A2 _04488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13535__I _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09674_ channels.atk_dec1\[7\] _01901_ _01905_ _02058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_94_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08877__A1 _01337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08625_ _01123_ _00029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10684__A1 _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08556_ _01071_ _01072_ _01073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10894__I _01104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08487_ net12 _01017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_49_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_162_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09108_ _01460_ _01560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_66_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10380_ _02522_ _02641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_60_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09039_ _01497_ _01498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12050_ clk_ctr\[0\] _02354_ _03732_ _00481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_92_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15925__I _07806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11001_ _03225_ _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_99_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12900__A3 _04905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10911__A2 _03052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09109__A2 _01560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14102__A2 _06055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13310__B1 _04784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15740_ _06291_ _07652_ _07655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08868__A1 channels.freq3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12952_ _04701_ _04707_ _04716_ _04958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_176_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13861__A1 _03284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11903_ _03905_ _03907_ _03985_ _03882_ _03986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_59_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10675__A1 channels.sample3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16756__I _00867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15671_ _03239_ _03237_ _07601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12883_ _03272_ _04242_ _04824_ _04889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_34_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15602__A2 _07529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17410_ _00480_ clknet_leaf_147_clk channels.adsr_state\[3\]\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14622_ _06527_ _06615_ _06616_ _06617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11834_ channels.env_counter\[0\]\[14\] channels.env_counter\[1\]\[14\] channels.env_counter\[2\]\[14\]
+ channels.env_counter\[3\]\[14\] _03886_ _01170_ _03925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_157_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17341_ _00411_ clknet_leaf_102_clk channels.freq2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11765_ _03834_ _03844_ _03855_ _03856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_3_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14553_ _06543_ _06548_ _06549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_99_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13180__I _05185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13504_ _04850_ _05510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10716_ _02936_ _02972_ _02973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_55_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14169__A2 _06062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17272_ _00342_ clknet_leaf_187_clk channels.accum\[2\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11696_ _03757_ _03781_ _03786_ _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14484_ _06355_ _06357_ _06481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_99_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_181_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_126_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16223_ _07727_ _08096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13435_ _05440_ _05281_ _05372_ _05441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10647_ _02900_ _02903_ _02905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10309__I channels.ch3_env\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer4 _04409_ net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_77_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16154_ spi_dac_i.spi_dat_buff_1\[5\] _07729_ _07921_ spi_dac_i.spi_dat_buff_1\[6\]
+ _03734_ _08030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_134_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_114_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13366_ _05369_ _05371_ _05372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_77_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10578_ _02792_ _02828_ _02836_ _02837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15669__A2 _07592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16866__A1 _03544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15105_ _07071_ _07072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_12317_ filters.cutoff_lut\[8\] filters.res_lut\[8\] _04217_ _04323_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_16085_ _07959_ _07962_ _07963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13297_ _05300_ _05301_ _05302_ _05303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_107_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_110_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12248_ _04253_ _04254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_15036_ _06980_ _07005_ _06979_ _00562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15835__I _07721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16618__A1 _01632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12179_ _04184_ _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09833__I _01750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16987_ _00066_ clknet_leaf_146_clk channels.accum\[0\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15841__A2 _07726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15938_ _07819_ _07820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13852__A1 _03284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10666__A1 _02505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15869_ _07750_ _07751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_149_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10130__A3 channels.pw3\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17608_ _00678_ clknet_leaf_168_clk _00010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09390_ _01788_ _01789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_149_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_3603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_164_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17539_ _00609_ clknet_leaf_201_clk channels.exp_periods\[3\]\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14186__I _01821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09587__A2 _01891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16857__A1 _02707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12343__A1 _04252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16609__A1 _01598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_35_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09743__I _01766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09726_ net11 _02098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09511__A2 _01899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09657_ channels.ctrl_reg2\[6\] _01974_ _01966_ channels.atk_dec2\[6\] _02041_ _02042_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_167_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08608_ channels.lfsr\[3\]\[8\] _01115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09588_ channels.freq3\[3\] _01870_ _01879_ channels.freq2\[3\] _01976_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08539_ _01019_ _01059_ _01025_ _01060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12609__I _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11550_ channels.freq2\[4\] _03670_ _03671_ _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_13_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11082__A1 filters.low\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_146_Left_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10501_ _02747_ _02754_ _02761_ _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_64_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09027__A1 _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11481_ _00389_ _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14020__A1 _06004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13220_ _05160_ _05161_ _05226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_107_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10432_ _02688_ _02690_ _02692_ _02693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_33_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12582__A1 _04574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17059__D _00129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16848__A1 _08419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13151_ _04165_ _04896_ _05155_ _05156_ _05157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_60_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10363_ _02623_ _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_103_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12102_ _03554_ channels.adsr_state\[1\]\[1\] _04131_ _04133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_20_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13082_ _05080_ _05081_ _05088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__14323__A2 _05487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10294_ _02554_ _02555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_72_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_1296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12334__A1 _04291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12033_ _04047_ _04090_ _04092_ _00472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16910_ _00984_ _00850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_155_Left_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12885__A2 _04890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16841_ tt_um_rejunity_sn76489.clk_counter\[2\] _00931_ _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10896__A1 _02366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14087__A1 _04645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16772_ _00884_ _00885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09189__S1 _01155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13984_ _05940_ _05956_ _05985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_176_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15723_ _07639_ _07643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12935_ _04287_ _04759_ _04941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_107_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15654_ _07498_ _07585_ _00600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_34_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12866_ _04772_ _04773_ _04872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_87_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14605_ _03396_ _06067_ _06600_ _06601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_11817_ _03905_ _03907_ _03908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__12519__I _04266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15585_ _07486_ _07520_ _07521_ _07522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_164_Left_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13062__A2 _04219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12797_ _04783_ _04803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_103_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17324_ _00394_ clknet_leaf_88_clk channels.freq1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14536_ _06527_ _06530_ _06531_ _06532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_11748_ _03828_ _03838_ _03839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16991__CLK clknet_5_28__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17255_ _00325_ clknet_leaf_76_clk filters.cutoff_lut\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09018__A1 channels.freq2\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09018__B2 channels.freq1\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14011__A1 _05512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14467_ _06462_ _06463_ _06464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11679_ channels.sus_rel2\[6\] _01280_ _01294_ channels.sus_rel1\[6\] _03770_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_55_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16206_ _07940_ _07820_ _08079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_154_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13418_ _05289_ _05377_ _05424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17186_ _00256_ clknet_leaf_105_clk channels.sus_rel3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_24_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14398_ net51 _06395_ _06396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XPHY_EDGE_ROW_180_Right_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12573__A1 _03302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10179__A3 channels.pw3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_5__f_clk_I clknet_3_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16137_ _07940_ _08011_ _08012_ _07912_ _08013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_45_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13349_ _05346_ _05354_ _05355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_3_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_149_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16068_ _07943_ _07946_ _07947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_173_Left_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_121_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_149_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15019_ _06987_ _06988_ _06989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_166_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08890_ _01257_ _01360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_166_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13085__I _04927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_127_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09511_ channels.sus_rel1\[0\] _01899_ _01901_ channels.atk_dec1\[0\] _01902_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_177_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_182_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09442_ _01825_ _01828_ _01832_ _01833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_78_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_182_Left_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_140_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09373_ _01773_ _01749_ _01763_ _01774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13053__A2 _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_163_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_31_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_160_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15502__A1 filters.mode_vol\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14305__A2 _06277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11119__A2 _03337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14069__A1 _06065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11508__I _03641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10342__A3 _02602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09709_ channels.freq1\[14\] _02082_ _02084_ _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_173_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10981_ _03201_ _03205_ _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__14819__I _05546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15018__B1 channels.sample2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12720_ _04457_ _04724_ _04725_ _04726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_167_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09422__B _01809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12651_ _04614_ _04656_ _04657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_66_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11602_ channels.pw3\[5\] _03704_ _03705_ _03707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_65_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12582_ _04574_ _04585_ _04588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_15370_ _07312_ _07322_ _07323_ _00578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_108_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14321_ _06317_ _06318_ _06319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11533_ _03657_ _03659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08471__A2 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17040_ _00110_ clknet_leaf_222_clk channels.lfsr\[1\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14252_ _06233_ _06250_ _06251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11464_ _01219_ _03616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10415_ _02644_ _02676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13203_ _04369_ _04882_ _05208_ _04320_ _05209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_11395_ channels.accum\[2\]\[12\] _03575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14183_ _06074_ _06181_ _06182_ _05869_ _06071_ _06183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_150_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10346_ _02503_ _02607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13134_ _05105_ _05108_ _05140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_104_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09971__A2 _02266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13065_ _05068_ _05070_ _05071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_40_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10277_ _02372_ _02538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_178_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09383__I net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12016_ channels.env_counter\[1\]\[2\] _04079_ _04082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_174_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_144_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16824_ _01776_ _00915_ _00921_ _00919_ _00827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_144_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13807__A1 _05792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_161_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_161_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16755_ _08449_ _00868_ _00872_ _00807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_105_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09487__A1 channels.ch3_env\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13967_ filters.low\[4\] _05969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_105_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15706_ _03216_ _03729_ _07628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_17_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12918_ _04923_ _04924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_85_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16686_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[7\] _08400_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[7\]
+ _08428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_122_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13898_ _05811_ _05900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_85_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15637_ _07562_ _07557_ _07569_ _07570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__12249__I _04254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12849_ _03364_ _04219_ _04854_ _04855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_146_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15568_ _07505_ _07506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_51_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17307_ _00377_ clknet_leaf_164_clk channels.accum\[1\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14519_ _06406_ _06513_ _06514_ _06515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_86_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15499_ _07438_ _07440_ _06913_ _07442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_141_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17238_ _00308_ clknet_leaf_13_clk filters.sample_filtered\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14535__A2 _04667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_168_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17169_ _00239_ clknet_leaf_145_clk channels.ctrl_reg3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_101_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09991_ _02234_ _02282_ _02285_ _00237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_122_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08942_ _01322_ _01406_ _01407_ _00062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12849__A2 _04219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_181_3735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_3746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09714__A2 _01891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08873_ _01338_ _01332_ _01343_ _01344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_93_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_179_3697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09425_ _01816_ _01817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14223__A1 _04326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09356_ filters.filt_2 _01758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14774__A2 _06761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09287_ _01712_ _01713_ _01706_ _01714_ _01145_ _01328_ _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_34_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09402__A1 _01767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10200_ _01582_ _02455_ channels.pw3\[0\] _02461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_28_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11180_ _03221_ _03395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_31_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10131_ _02390_ channels.pw2\[11\] _01096_ _02392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_101_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10062_ _02308_ _02331_ _02336_ _00257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09261__S0 _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14870_ _06849_ _06850_ _00551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13821_ _05819_ _05823_ _05824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_173_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09469__A1 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14462__A1 _04576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16540_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[0\] _08322_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[0\]
+ _08323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_67_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13752_ _05644_ _05645_ _05649_ _05756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10964_ filters.filter_step\[2\] _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_70_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12703_ _04265_ _04491_ _04709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12069__I _04106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16471_ _08262_ _08264_ _07740_ _00738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13683_ _05588_ _05687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14214__A1 _04896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10895_ channels.sample2\[0\] _03143_ _03144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15422_ _06837_ _07365_ _07362_ _07370_ _07371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_12634_ _04628_ _04631_ _04636_ _04638_ _04640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_182_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12776__A1 _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15353_ _07306_ _07300_ _07307_ _07308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_136_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09641__A1 channels.pw1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12565_ _04297_ _04498_ _04571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09641__B2 channels.ctrl_reg1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14304_ _06281_ _06301_ _06299_ _06173_ _06302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_163_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11516_ _03513_ _03642_ _03647_ _00400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_124_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15284_ _07227_ _07230_ _07244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_12496_ _04499_ _04501_ _04502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_145_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17023_ _00000_ clknet_leaf_240_clk filters.res_lut\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10317__I channels.ch3_env\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14235_ _06128_ _06132_ _06234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_151_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12733__S _04710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11447_ channels.accum\[1\]\[9\] _03605_ _03606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_180_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_1263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11200__A1 _03411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14166_ _05979_ _06058_ _06166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_46_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11378_ _03138_ _01381_ _03564_ _00345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13117_ _03349_ _04315_ _04191_ _05123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10329_ _02589_ _02590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14097_ _04416_ _06096_ _06097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_163_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16690__A2 _08289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13048_ _04946_ _05054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12700__A1 _04705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08904__B1 _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10052__I _01818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16807_ _01756_ _00906_ _00909_ _00910_ _00821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_1_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17787_ _00857_ clknet_leaf_56_clk tt_um_rejunity_sn76489.control_noise\[0\]\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_163_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14999_ _06939_ _05035_ _05040_ _06970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_16738_ _08463_ _00861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09062__B _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16669_ _08413_ _08414_ _00786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09880__A1 _02160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09210_ _01647_ _01648_ _01639_ _01649_ _01643_ _01644_ _01650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_8_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17685__CLK clknet_5_11__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09141_ _01043_ _01588_ _01590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_29_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12707__I _04712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11611__I _03711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09072_ _01527_ _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_47_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_135_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09935__A2 _01833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09974_ _02270_ _02265_ _02271_ _02273_ _00232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_110_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08925_ _01391_ _01392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09699__A1 _01767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08856_ _01158_ _01328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__13247__A2 _04712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14444__A1 _04318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08787_ channels.accum\[0\]\[0\] _01260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13273__I _05077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09408_ _01792_ _01803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10680_ _02895_ _02926_ _02928_ _02937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_165_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09339_ _01741_ _01742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09623__A1 channels.ch3_env\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_109_Right_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_152_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09623__B2 channels.atk_dec1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12350_ _04354_ _04355_ _04356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_69_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11430__B2 _03592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11301_ _02316_ _03498_ _03504_ _00328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_12281_ _04286_ _04287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_50_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14020_ _06004_ _06020_ _06021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__13183__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11232_ _03235_ _03442_ _03443_ _03444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_31_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12930__A1 _04632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11163_ _03283_ _03379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_8_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10114_ channels.ctrl_reg1\[2\] channels.ring_outs\[2\] _01284_ _02375_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_101_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15971_ _07795_ _07786_ _07851_ _07852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11094_ filters.band\[5\] _03314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_179_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17710_ _00780_ clknet_leaf_232_clk channels.lfsr\[0\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10045_ _02319_ _02320_ _02323_ _00253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11497__A1 channels.freq1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14922_ _05547_ _06897_ _06898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_141_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17641_ _00711_ clknet_leaf_204_clk channels.ch3_env\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_76_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14853_ _06799_ _06831_ _06832_ _06752_ _06834_ _06835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_26_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14435__A1 _06417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13804_ _05804_ _05805_ _05806_ _05807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__11249__A1 _03236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17572_ _00642_ clknet_5_5__leaf_clk filters.filter_step\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_98_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14986__A2 _06949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14784_ _06754_ _06772_ _06773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11996_ _03900_ _03911_ _04058_ _04066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_86_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_82_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16523_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[8\] _08270_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[8\]
+ _08309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_82_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13735_ _05717_ _05738_ _05739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10947_ _03174_ _03104_ _03175_ _00303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09862__A1 _02179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16454_ _07683_ _08252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_156_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13666_ _04500_ _05663_ _05670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14738__A2 _06397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_205_clk_I clknet_5_23__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10878_ _03112_ _03115_ _03129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_144_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_94_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15405_ _07355_ _07356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12617_ _04614_ _04621_ _04622_ _04623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_16385_ _08196_ _08199_ _08200_ _00716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_156_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13597_ _05582_ _05601_ _05602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_53_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13410__A2 _05415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15336_ filters.low\[18\] _06396_ _07292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_81_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12548_ _04551_ _04553_ _04554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_117_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15267_ _07210_ _07215_ _07228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_2 _01588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12479_ _04267_ _04485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_22_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17006_ _00085_ clknet_leaf_224_clk channels.lfsr\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13174__A1 filters.band\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14218_ _06129_ _06130_ _06217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_1_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15198_ _07152_ _07156_ _07161_ _07162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_0_111_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14149_ _06015_ _06016_ _06149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_6_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_130_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09225__S0 _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08710_ _01176_ channels.exp_periods\[3\]\[4\] _01194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11488__A1 channels.freq1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09690_ _01781_ _01970_ _02073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_83_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08641_ _01131_ _00037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer14 _06709_ net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10160__A1 _01555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer25 net65 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__10160__B2 _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer36 _06835_ net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_179_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14977__A2 _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08572_ _01088_ _01089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12988__A1 _04512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11335__S1 _01160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_176_3645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09853__A1 channels.pw2\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_176_3656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12452__A3 _04376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09124_ channels.lfsr\[0\]\[17\] _01573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_40_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09081__A2 _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16353__B _01821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09055_ _01504_ _01502_ _01511_ _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__16351__A1 _02356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15154__A2 _07119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12212__I0 filters.cutoff_lut\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12912__A1 _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_38_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09957_ _02240_ _02257_ _02261_ _00227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08908_ channels.freq2\[5\] _01276_ _01288_ channels.freq1\[5\] _01376_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_09888_ _02185_ _02210_ _02213_ _00206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_99_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08839_ _01308_ channels.accum\[3\]\[0\] _01312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10151__A1 channels.pw1\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11850_ _03744_ _03937_ _03940_ _03941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_135_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16528__B _08313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10801_ _03049_ _03050_ _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_95_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09844__A1 channels.pw2\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11781_ _03804_ _03825_ _03872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13520_ _05456_ _05459_ _05525_ _05526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_83_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10454__A2 _02710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10732_ _02952_ _02958_ _02988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13451_ _05303_ _05332_ _05457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_48_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10663_ _01715_ _02771_ _02921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12402_ _04398_ _04399_ _04407_ _04408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_16170_ _08017_ _08021_ _08045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_51_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11403__A1 _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13382_ _04941_ _05386_ _05387_ _05388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10594_ _02575_ _02589_ _02853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_191_clk_I clknet_5_22__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15121_ _07082_ _07085_ _07087_ _07088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_106_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12333_ _04331_ _04338_ _04339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_23_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_3_0_clk clknet_0_clk clknet_3_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_clkbuf_leaf_71_clk_I clknet_5_14__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15052_ _07018_ _07019_ _07020_ _07021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_105_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12264_ _04266_ _04269_ _04270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14003_ _05908_ _05917_ _06003_ _06004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_31_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11200__B _03413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11215_ _03427_ _03428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_112_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12195_ _04200_ _04201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_75_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_75_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_112_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11146_ _03362_ _03363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_clkbuf_leaf_86_clk_I clknet_5_12__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15954_ _07834_ _07835_ _07836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11077_ filters.high\[4\] _03298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_10028_ _02309_ _02311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14905_ filters.low\[29\] _06882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_15885_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[3\] _07766_ _07767_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__14408__A1 _06373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_196_clk clknet_5_23__leaf_clk clknet_leaf_196_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10142__A1 _01085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10142__B2 _02402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11426__I _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17624_ _00694_ clknet_leaf_209_clk channels.env_vol\[1\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14836_ _06760_ _06820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_1254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_158_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17555_ _00625_ clknet_leaf_23_clk filters.low\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14767_ _06754_ _06756_ _06757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_11979_ _04043_ _04051_ _04052_ _00458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_144_clk_I clknet_5_30__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16506_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[5\] _08269_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[5\]
+ _08295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_85_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11642__A1 channels.clk_div\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13718_ _03383_ _04342_ _05721_ _05722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_128_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08735__I _01100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17486_ _00556_ clknet_leaf_27_clk filters.band\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_160_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14698_ _06599_ _06601_ _06693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_119_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_154_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16437_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[0\] _08238_ _08239_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_27_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13649_ _03251_ _05545_ _05652_ _05653_ _00527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__11161__I _03376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_171_3553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_171_3564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16368_ _03974_ _08184_ _08187_ _00712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_159_clk_I clknet_5_28__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15319_ _07270_ _07272_ _07273_ _07276_ _07277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_169_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16299_ channels.env_counter\[3\]\[5\] _08147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_140_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_132_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_39_clk_I clknet_5_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09811_ _02157_ _02151_ _02159_ _00183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08574__B2 channels.ring_outs\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16399__I _08194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09742_ _02110_ _02107_ _02111_ _00162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_158_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09673_ channels.ctrl_reg2\[7\] _01830_ _01904_ _02056_ _02057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_187_clk clknet_5_19__leaf_clk clknet_leaf_187_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11336__I _03529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13870__A2 _05657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08624_ channels.lfsr\[3\]\[16\] _01123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10240__I _02500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08555_ channels.clk_div\[1\] _01072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09826__A1 _02131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13622__A2 _05624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_59_Left_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08486_ _01015_ _01016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_147_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_175_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15375__A2 _06599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09107_ _01323_ _01557_ _01558_ _01559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_32_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14382__I filters.band\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_111_clk clknet_5_15__leaf_clk clknet_leaf_111_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09476__I _01866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09038_ channels.accum\[0\]\[14\] channels.accum\[1\]\[14\] channels.accum\[2\]\[14\]
+ channels.accum\[3\]\[14\] _01495_ _01496_ _01497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_131_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_68_Left_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_131_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_92_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11000_ _03224_ _03225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_99_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10372__A1 _01305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_70_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12951_ _04456_ _04460_ _04957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_leaf_178_clk clknet_5_18__leaf_clk clknet_leaf_178_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_99_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11902_ _03983_ _03921_ _03984_ _03985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_15670_ _07599_ _07595_ _07600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12882_ _03287_ _04196_ _04803_ _04888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_158_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_77_Left_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_14621_ _06356_ _06473_ _06530_ _06616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11833_ _03850_ _03814_ _03890_ _03924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_96_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17340_ _00410_ clknet_leaf_100_clk channels.freq2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14552_ _06546_ _06547_ _06548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11764_ _03853_ _03854_ _03855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_161_Right_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_99_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13503_ _04848_ _05509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10715_ _02937_ _02971_ _02972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_17271_ _00341_ clknet_leaf_178_clk channels.accum\[2\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__16772__I _00884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14483_ _06380_ _05563_ _06480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11695_ channels.atk_dec3\[0\] _03782_ _03783_ channels.atk_dec2\[0\] _03785_ _03786_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_148_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16222_ _07726_ _08094_ _08095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_64_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13434_ _04562_ _05440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10646_ _02900_ _02903_ _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_181_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16153_ _08007_ _08026_ _08028_ _08029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_141_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer5 _04346_ net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_114_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_102_clk clknet_5_13__leaf_clk clknet_leaf_102_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_114_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13365_ _04641_ _05370_ _05371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_77_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10577_ _02794_ _02827_ _02836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_77_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15104_ _07045_ _07046_ _07070_ _07071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12316_ _04321_ _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16084_ _07960_ _07961_ _07781_ _07962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16866__A2 _03755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13296_ _05207_ _05225_ _05302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15035_ _06983_ _07004_ _07005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12247_ _04235_ _04253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_43_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12178_ filters.res_lut\[0\] _04167_ _04184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_78_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11129_ filters.band\[7\] _03347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_16986_ _00065_ clknet_leaf_152_clk channels.accum\[0\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15937_ _07817_ _07818_ _07819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_169_clk clknet_5_24__leaf_clk clknet_leaf_169_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_79_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10060__I _02334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15868_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[1\] _07745_ _07750_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10666__A2 _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17607_ _00677_ clknet_leaf_162_clk _00009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14819_ _05546_ _06804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_148_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15799_ _07663_ _07698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14801__A1 _06706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11615__A1 channels.pw2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17538_ _00608_ clknet_leaf_202_clk channels.exp_periods\[3\]\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_171_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17469_ _00539_ clknet_leaf_15_clk filters.band\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09296__I _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08547__A1 clk_trg\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_5_28__f_clk clknet_3_7_0_clk clknet_5_28__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_10_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_35_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09725_ channels.pw1\[11\] _02097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_5_22__f_clk_I clknet_3_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15761__I _07639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09656_ _01908_ _02038_ _02039_ _02040_ _02041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_69_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08607_ _01114_ _00020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_167_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09587_ channels.pw1\[11\] _01891_ _01975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08538_ _01036_ _01044_ _01059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_182_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08469_ net6 _00998_ _00999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_9_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13359__A1 _04420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10500_ _02755_ _02760_ _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11480_ _03623_ _00389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10431_ _02667_ _02668_ _02691_ _02692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_94_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12625__I _04630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13150_ _05111_ _05112_ _05156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_143_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10362_ _02622_ _02623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_60_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12101_ _04132_ _00500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13081_ _04288_ _05049_ _05087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10293_ _02553_ _02554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_72_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09934__I _02104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12334__A2 _04266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12032_ channels.env_counter\[1\]\[8\] _04091_ _04092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12360__I _04323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16840_ _06917_ _00930_ _00931_ _00833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__10896__A2 _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15284__A1 _07227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16771_ _00879_ _00883_ _00884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13983_ _05981_ _05983_ _05984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_137_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15722_ _05759_ _07637_ _07642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12934_ _04844_ _04868_ _04939_ _04940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_107_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_107_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15653_ filters.sample_buff\[10\] _07447_ _07523_ _07584_ _07585_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_12865_ _04814_ _04870_ _04871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14604_ filters.low\[10\] _03377_ _06600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11816_ _03906_ _03816_ _03836_ _03907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_68_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15584_ _07512_ _07507_ _07519_ _07521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_29_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12796_ _04801_ _04802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_157_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13062__A3 _04403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17323_ _00393_ clknet_leaf_77_clk channels.freq1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_28_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14535_ _06356_ _04667_ _06531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11747_ _03802_ _03813_ _03838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17254_ _00324_ clknet_leaf_75_clk filters.cutoff_lut\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_14466_ _05510_ _05989_ _06463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11678_ channels.sus_rel3\[6\] _01081_ _03769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16205_ _07983_ _07749_ _08078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13417_ _05037_ _05043_ _05048_ _05422_ _05423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_70_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17185_ _00255_ clknet_leaf_105_clk channels.sus_rel3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10629_ _02842_ _02877_ _02887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_180_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_14397_ _06390_ _06394_ _06395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_16136_ _07825_ _07906_ _08012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13770__A1 _04630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12573__A2 _04332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13348_ _05348_ _05353_ _05354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_51_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16451__B _08098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16067_ _07880_ _07944_ _07945_ _07946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_11_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13279_ _05271_ _05274_ _05284_ _05285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_149_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15018_ _01744_ channels.sample1\[3\] channels.sample2\[3\] _01758_ _06988_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_166_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_166_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10887__A2 _03136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16969_ _00048_ clknet_leaf_191_clk channels.exp_counter\[1\]\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09510_ _01900_ _01901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14873__I1 _06472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15027__A1 filters.low\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09441_ _01831_ _01832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_182_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_140_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09372_ _01772_ _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_75_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12261__A1 _03348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12445__I _04450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15502__A2 _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13513__A1 _04850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10590__A4 _02847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10327__A1 _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12180__I _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08940__A1 _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15491__I _06978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09708_ _01807_ _02081_ _02085_ _00154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10980_ _03202_ _03204_ _03205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_97_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09639_ channels.freq3\[5\] _01937_ _01999_ channels.ctrl_reg3\[5\] _02025_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_97_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12650_ _04644_ _04620_ _04618_ _04656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11601_ _03668_ _03703_ _03706_ _00426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_66_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12581_ _04559_ _04560_ _04586_ _04587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_93_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_14320_ _06207_ _06208_ _06318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_66_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11532_ _03657_ _03658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08833__I _01305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14251_ _06236_ _06249_ _06250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_80_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11463_ _01104_ _03615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_151_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13202_ _05107_ _05208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10414_ _02599_ _02514_ _02662_ _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_1_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14182_ _05972_ _06070_ _06071_ _06182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_11394_ _03566_ _01459_ _03574_ _00351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13133_ _04369_ _04818_ _05139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10345_ _02597_ _02605_ _02606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13064_ _03382_ _05069_ _04341_ _05070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_10276_ _02524_ _02528_ _02536_ _02537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XPHY_EDGE_ROW_70_Right_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12015_ _04017_ _04076_ _04081_ _00465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_5_11__f_clk clknet_3_2_0_clk clknet_5_11__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_109_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16823_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[3\] _00916_ _00921_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_144_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_161_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16754_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[5\] _00869_ _00871_ _00872_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13966_ _05877_ _05967_ _05968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_45_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12917_ _04861_ _04923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15705_ _07627_ _00609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16685_ _08419_ _08427_ _00789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_122_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13897_ _05886_ _05898_ _05899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_85_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15636_ filters.sample_buff\[9\] _07568_ _07569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12848_ _04271_ _04854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09239__A2 _01659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14232__A2 _06155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15567_ filters.sample_buff\[4\] _07504_ _07505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_14_Left_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12779_ _03253_ _04225_ _04784_ _04785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_56_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17306_ _00376_ clknet_leaf_152_clk channels.accum\[1\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14518_ _06409_ _06489_ _06514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_12_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15498_ _07438_ _07440_ _07441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_28_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14449_ _06432_ _06445_ _06446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_17237_ _00307_ clknet_5_6__leaf_clk filters.sample_filtered\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_154_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15732__A2 _07632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13743__A1 _05743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17168_ _00238_ clknet_leaf_145_clk channels.ctrl_reg3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_168_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16119_ _07994_ _07995_ _07996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_12_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17099_ _00169_ clknet_leaf_111_clk channels.atk_dec1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09990_ channels.ctrl_reg3\[4\] _02283_ _02284_ _02285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08941_ channels.accum\[0\]\[7\] _01360_ _01407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_181_3736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08872_ _01341_ _01342_ _01343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_181_3747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_91_clk clknet_5_7__leaf_clk clknet_leaf_91_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09424_ net15 _01816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_48_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_179_3698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09355_ _01756_ _01757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_47_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09749__I _02106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13982__A1 _05982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09286_ channels.lfsr\[3\]\[20\] _01714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09484__I _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_1197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10130_ _02389_ _02390_ channels.pw3\[11\] _02391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_30_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11519__I _03641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10061_ filters.cutoff_lut\[9\] _02332_ _02335_ _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_89_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09261__S1 _01680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08913__A1 _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13820_ _05820_ _05821_ _05822_ _05823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_3_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14462__A2 _05990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13751_ _05754_ _05755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10963_ _03187_ _03188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_98_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_82_clk clknet_5_9__leaf_clk clknet_leaf_82_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_134_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12702_ _04701_ _04707_ _04708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16470_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[0\] _08263_ _08264_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13682_ _05607_ _05615_ _05685_ _05686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_10894_ _01104_ _03143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14214__A2 _05181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15421_ _07365_ _07364_ _07370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_182_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12633_ _04628_ _04631_ _04636_ _04638_ _04639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XTAP_TAPCELL_ROW_100_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13422__B1 _05417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10236__B1 channels.ctrl_reg1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15352_ _07295_ _06294_ _07292_ _07307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_80_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12564_ _04564_ _04568_ _04569_ _04570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_80_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14303_ _06275_ _06277_ _06301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_109_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11515_ channels.pw1\[2\] _03643_ _03644_ _03647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15283_ _07242_ _07243_ _00571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__15714__A2 _03730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12495_ _04301_ _04500_ _04425_ _04501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_163_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17022_ _00101_ clknet_leaf_212_clk channels.lfsr\[2\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13725__A1 _04274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14234_ _06231_ _06232_ _06233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12528__A2 _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11446_ _03149_ _03605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12813__I _04818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14165_ _05979_ _06058_ _06165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11377_ channels.accum\[2\]\[5\] _03559_ _03564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13116_ _04367_ _04290_ _05122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10328_ _02484_ _02498_ _02588_ _02589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_81_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14096_ _06005_ _06096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_163_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13047_ _04643_ _05049_ _05052_ _05053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10333__I _02544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10259_ channels.env_vol\[0\]\[2\] channels.env_vol\[1\]\[2\] _02519_ _02520_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_56_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16806_ _02102_ _00910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17786_ _00856_ clknet_leaf_205_clk channels.exp_periods\[0\]\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14998_ filters.low\[3\] _06968_ _06969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_152_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16737_ _08449_ _08464_ _00860_ _00801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_163_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13949_ _04229_ _05351_ _05951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_73_clk clknet_5_14__leaf_clk clknet_leaf_73_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_147_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16668_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[3\] _08345_ _01753_ _08414_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Left_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15619_ channels.sample1\[8\] _03427_ _07553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16599_ _08356_ _08372_ _00758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09140_ _01588_ _01589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_84_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09632__A2 _02017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_139_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09071_ channels.accum\[0\]\[17\] channels.accum\[1\]\[17\] channels.accum\[2\]\[17\]
+ channels.accum\[3\]\[17\] _01139_ _01480_ _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_114_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13716__A1 _04802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_135_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_31_Left_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09973_ _02272_ _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11339__I _03532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10950__A1 channels.sample1\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10243__I _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08924_ _01389_ _01390_ _01391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_110_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08855_ _01325_ _01326_ _01327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_100_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08786_ _01259_ _00054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_93_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input13_I bus_in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12455__A1 _04456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_40_Left_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_64_clk clknet_5_11__leaf_clk clknet_leaf_64_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_138_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_45_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09407_ _01792_ _01802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14385__I _06261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09338_ _01740_ _01741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__13955__A1 _05940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09269_ channels.lfsr\[2\]\[18\] _01700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_30_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_161_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11300_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[2\] _03500_ _03503_ _03504_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12280_ filters.res_lut\[3\] _04169_ _04286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_105_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13183__A2 _05184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11231_ filters.high\[13\] _03235_ _03443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09428__B _01809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11162_ _03377_ _03378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_140_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10941__A1 channels.sample1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09139__A1 _01581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10113_ channels.ctrl_reg3\[2\] channels.ring_outs\[1\] _01073_ _02374_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_105_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15970_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[0\] _07788_ _07851_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11093_ _03195_ _03313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_175_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10044_ channels.sus_rel3\[4\] _02321_ _02322_ _02323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14921_ _06722_ _06893_ net70 _06897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__12694__A1 _04699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17640_ _00710_ clknet_leaf_207_clk channels.ch3_env\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_14852_ _06814_ _06816_ _06825_ _06833_ _06834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__14435__A2 _06431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13803_ _04221_ _05187_ _05806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17571_ _00641_ clknet_leaf_22_clk filters.low\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14783_ filters.low\[17\] filters.band\[17\] _06755_ _06772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11995_ _04007_ _04064_ _04065_ _00461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_55_clk clknet_5_8__leaf_clk clknet_leaf_55_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_82_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16522_ _08307_ _08308_ _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13734_ _05719_ _05737_ _05738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__12997__A2 _05000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10946_ channels.sample1\[8\] _03170_ _03175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16453_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[4\] _08249_ _08251_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_27_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13665_ _05667_ _05668_ _05669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_39_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10877_ _03031_ _03128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_155_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15404_ _02100_ _07355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12749__A2 _04743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13946__A1 _04238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12616_ _04541_ _04618_ _04622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16384_ _08195_ _08200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13946__B2 _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09075__B1 _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_156_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13596_ _05584_ _05600_ _05601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_26_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15335_ filters.low\[17\] _06293_ _07291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12547_ _04352_ _04359_ _04552_ _04553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_108_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15266_ _07212_ _07213_ _07226_ _07227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_12478_ _04174_ _04483_ _04484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_3 _01590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09378__A1 filters.res_filt\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11709__C2 channels.atk_dec1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17005_ _00084_ clknet_leaf_219_clk channels.lfsr\[2\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14217_ _06201_ _06215_ _06216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13174__A2 _05179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11429_ channels.accum\[1\]\[2\] _03595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_112_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15197_ _07157_ _07160_ _07161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_158_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_9__f_clk clknet_3_2_0_clk clknet_5_9__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14148_ _06015_ _06016_ _06148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_21_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_130_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14079_ _03314_ _05545_ _06079_ _05653_ _00531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09225__S1 _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input5_I addr[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08640_ channels.env_vol\[3\]\[1\] _01131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_175_Right_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08468__I net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14426__A2 _05075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer15 _05375_ net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer26 _05378_ net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__15803__B _07700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer37 _05413_ net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__12437__A1 filters.cutoff_lut\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08571_ _01087_ _01083_ _01088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_17769_ _00839_ clknet_leaf_203_clk channels.exp_periods\[2\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_46_clk clknet_5_2__leaf_clk clknet_leaf_46_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_53_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12988__A2 _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_159_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_176_3646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_176_3657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11622__I _03711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09161__S0 _01605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09123_ _01540_ _01571_ _01572_ _00078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_162_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09081__A3 _01534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09054_ _01504_ _01502_ _01511_ _01512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_115_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10923__A1 channels.sample2\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09956_ channels.freq3\[14\] _02258_ _02255_ _02261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15862__A1 _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08907_ channels.freq3\[5\] _01076_ _01375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09887_ channels.atk_dec2\[1\] _02211_ _02206_ _02213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09541__A1 _01823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08838_ channels.accum\[2\]\[0\] _01311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_142_Right_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_135_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_174_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08769_ _01088_ _01245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14968__A3 channels.sample1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_37_clk clknet_5_3__leaf_clk clknet_leaf_37_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_67_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10800_ _02358_ _03054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11780_ _03824_ _03870_ _03871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10731_ _02960_ _02966_ _02964_ _02987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_177_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12628__I _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13450_ _05442_ _05455_ _05456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_94_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10662_ _02402_ _02567_ _02920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_125_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12401_ _04401_ _04406_ _04407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13381_ _04643_ _05054_ _04944_ _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_134_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10593_ _02508_ _02513_ _02637_ _02852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_23_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15120_ _07082_ _07085_ _07086_ _07087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_106_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12332_ _04334_ _04337_ _04338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_63_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13459__I _05229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15051_ _01746_ channels.sample1\[4\] _07020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12263_ _04268_ _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_160_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14002_ _05912_ _05916_ _06003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11214_ _03401_ _03427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12194_ _04199_ _04200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_82_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11145_ _03191_ _03248_ _03197_ _03361_ _03362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XANTENNA__09672__I channels.sample3\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15953_ _07764_ _07832_ _07835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_37_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11076_ filters.sample_filtered\[4\] _03297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_179_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09532__A1 channels.pw1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10027_ _02309_ _02310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09532__B2 channels.freq1\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14904_ _06880_ _06881_ _00554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_15884_ _07765_ _07766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_153_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17623_ _00693_ clknet_leaf_128_clk channels.env_counter\[3\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14835_ _06804_ _06818_ _06819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11890__A2 _03974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_158_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17554_ _00624_ clknet_leaf_25_clk filters.low\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_158_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11978_ channels.env_counter\[2\]\[9\] _04048_ _04052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14766_ filters.low\[16\] filters.band\[16\] _06755_ _06756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16505_ _08265_ _08294_ _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13717_ _04825_ _05721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_50_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10929_ channels.sample1\[1\] _03164_ _03165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_168_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17485_ _00555_ clknet_leaf_246_clk filters.band\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14697_ _06689_ _06691_ _06692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_156_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_119_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_156_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16436_ _08237_ _08238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13648_ _01822_ _05653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_171_3554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10058__I _01750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13579_ _05464_ _05474_ _05583_ _05584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_16367_ channels.ch3_env\[5\] _08185_ _08187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_171_3565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09847__I _02184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15318_ _07274_ _07264_ _07275_ _07276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_16298_ _08146_ _00683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_124_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08810__A3 _01282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_132_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13147__A2 _05124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_10_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12273__I _04278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15249_ _01772_ channels.sample3\[11\] _07211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_99_Right_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__16097__A1 _07838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09810_ channels.sus_rel1\[6\] _02152_ _02158_ _02159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08574__A2 _01086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15844__A1 _04776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09741_ channels.ctrl_reg1\[1\] _02108_ _02094_ _02111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09523__A1 filters.cutoff_lut\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09523__B2 filters.cutoff_lut\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09672_ channels.sample3\[11\] _02056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11330__A1 _03511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08623_ _01122_ _00028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13870__A3 _05849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_19_clk clknet_5_3__leaf_clk clknet_leaf_19_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10684__A3 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08554_ channels.clk_div\[2\] _01071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_49_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13083__A1 _05080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_6_Left_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11633__A2 _01093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10436__A3 _02686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08485_ _01010_ _01012_ _01014_ _01015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_92_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14583__A1 _04806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09106_ _01554_ _01556_ _01558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08661__I _01144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09037_ _01153_ _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12897__A1 _03316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_92_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11728__S _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_204_clk_I clknet_5_22__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09939_ _02245_ _02247_ _02249_ _00221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_70_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13310__A2 _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12950_ _04953_ _04954_ _04955_ _04956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_70_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11901_ _03923_ _03926_ _03984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_29_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12881_ _03302_ _04332_ _04800_ _04887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_clkbuf_leaf_219_clk_I clknet_5_21__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11832_ _03915_ _03920_ _03923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14620_ _06614_ _06473_ _06530_ _06615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13074__A1 _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14551_ _06544_ _06545_ _06547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11763_ channels.env_counter\[0\]\[6\] channels.env_counter\[1\]\[6\] channels.env_counter\[2\]\[6\]
+ channels.env_counter\[3\]\[6\] _03832_ _03842_ _03854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__10427__A3 _02687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13502_ _05502_ _05507_ _05508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10714_ _02942_ _02970_ _02971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_95_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_166_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14482_ _06477_ _06478_ _06479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17270_ _00340_ clknet_leaf_182_clk channels.accum\[2\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11694_ _03784_ _03785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_55_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16221_ _08077_ _08092_ _08094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13433_ _05436_ _05437_ _05438_ _05439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__14574__A1 _04893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10645_ _02901_ _02902_ _02903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_64_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16152_ _07987_ _08000_ _08027_ _08028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_106_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13364_ _05367_ _05370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_91_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10576_ _02788_ _02833_ _02834_ _02835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_63_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer6 _05423_ net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_77_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12315_ _04320_ _04321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15103_ _01770_ _01927_ _07047_ _07070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_16083_ _07890_ _07778_ _07961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_122_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13295_ _05240_ _05301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__16866__A3 _00953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15034_ _07001_ _07003_ _07004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12246_ _04244_ _04250_ _04251_ _04252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__12888__A1 _04893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09753__A1 channels.ctrl_reg1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12177_ _04176_ _04182_ _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11560__A1 _03677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15826__A1 _03735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11128_ _03218_ _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16985_ _00064_ clknet_leaf_163_clk channels.accum\[0\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15936_ tt_um_rejunity_sn76489.chan\[3\].attenuation.in _07818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_11059_ filters.sample_filtered\[3\] _03281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_155_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11312__A1 _03511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15867_ _07748_ _07749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17606_ _00676_ clknet_leaf_48_clk net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_176_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09351__B _01753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14818_ _06802_ _06803_ _00546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_114_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15798_ _07636_ _07697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_86_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17537_ _00607_ clknet_leaf_215_clk channels.exp_periods\[3\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14749_ _03468_ _06710_ _06740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17468_ _00538_ clknet_leaf_26_clk filters.band\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_15_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16419_ _08224_ _08225_ _08222_ _00725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_156_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14565__A1 _06417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17399_ _00469_ clknet_leaf_138_clk channels.env_counter\[1\]\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10051__A1 _02326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09992__A1 channels.ctrl_reg3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08795__A2 channels.ctrl_reg2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16857__A3 _03128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_8_clk clknet_5_5__leaf_clk clknet_leaf_8_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_140_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12731__I _04711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11551__A1 _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09724_ _01767_ _02090_ _02096_ _00159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11303__A1 _02299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10106__A2 _01560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09655_ channels.atk_dec3\[6\] _01991_ _01992_ channels.freq3\[14\] _02040_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_190_clk_I clknet_5_22__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08606_ channels.lfsr\[3\]\[7\] _01114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_3_2_0_clk clknet_0_clk clknet_3_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_09586_ _01829_ _01974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13056__A1 _04900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08656__I _01139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_70_clk_I clknet_5_14__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08537_ _01057_ _01058_ _00004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08468_ net5 _00998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__11015__C _03239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09680__B1 _01937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13359__A2 _05281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10290__A1 _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_85_clk_I clknet_5_12__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10430_ _02681_ _02682_ _02691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_61_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_94_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_94_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09983__A1 channels.ctrl_reg3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10426__I _02686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10361_ _02538_ _02619_ _02621_ _02499_ _02622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_61_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12100_ _03545_ channels.adsr_state\[1\]\[0\] _04131_ _04132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13080_ net41 _05084_ _05085_ _05086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10292_ _02484_ _02498_ _02552_ _02553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_103_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09735__A1 _01781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12031_ _04077_ _04091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_72_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_143_clk_I clknet_5_27__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11542__A1 _03664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_23_clk_I clknet_5_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15952__I _07726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15284__A2 _07230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16770_ _08441_ _08462_ _00880_ _00881_ _00882_ _00883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_13982_ _05982_ _05883_ _05896_ _05983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13834__A3 _05731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15721_ _07638_ _07641_ _00611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_158_clk_I clknet_5_28__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12933_ _04846_ _04867_ _04939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_77_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11845__A2 _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_107_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_38_clk_I clknet_5_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15652_ _07582_ _07583_ _07584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12864_ _04840_ _04869_ _04870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_69_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14603_ _06512_ _06598_ _06599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_96_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11815_ _03828_ _03906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15583_ _07512_ _07507_ _07519_ _07520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_12795_ _04800_ _04801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_69_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17322_ _00392_ clknet_leaf_77_clk channels.freq1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_55_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11746_ _03794_ _03837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14534_ _06454_ _06528_ _06529_ _06530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_172_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16536__A2 _08315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10281__A1 _01482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17253_ _00323_ clknet_leaf_75_clk filters.cutoff_lut\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_12_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14465_ _05509_ _05793_ _06462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11677_ _01168_ _02533_ _03767_ _03768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_16204_ _08069_ _08071_ _08076_ _08077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_114_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10628_ _02844_ _02876_ _02886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13416_ net55 _05404_ _05416_ _05421_ _05422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_109_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17184_ _00254_ clknet_leaf_104_clk channels.sus_rel3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_24_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14396_ _06391_ _06393_ _06394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_181_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10033__A1 channels.sus_rel3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16135_ _07825_ _07906_ _07846_ _08011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_148_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13347_ _05349_ _05352_ _05353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_51_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__16839__A3 _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10559_ _02817_ _02818_ _02819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__12573__A3 _04578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16066_ _07903_ _07914_ _07945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13278_ _05275_ _05283_ _05284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_80_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12229_ filters.cutoff_lut\[7\] filters.res_lut\[7\] _04217_ _04235_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15017_ filters.filt_2 filters.filt_1 channels.sample1\[3\] channels.sample2\[3\]
+ _06987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_TAPCELL_ROW_166_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13583__S _05179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10071__I _02334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_127_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16968_ _00047_ clknet_leaf_192_clk channels.exp_counter\[1\]\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_155_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_159_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15919_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[0\] _07801_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11836__A2 _03925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16899_ _00969_ channels.exp_periods\[1\]\[3\] _00975_ _00979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09440_ net4 net3 _01831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__13038__A1 _04952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09371_ _01771_ _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_176_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12261__A2 _04190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_96_Left_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_145_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_172_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10024__A1 _02242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09965__A1 _02245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09717__A1 channels.pw1\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12461__I _04254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14710__A1 _06703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11524__A1 _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10327__A2 _02381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09707_ channels.freq1\[13\] _02082_ _02084_ _02085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_69_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15018__A2 channels.sample1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09638_ channels.pw2\[5\] _01996_ _01997_ channels.freq2\[13\] _02024_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_139_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09569_ channels.atk_dec2\[2\] _01837_ _01895_ channels.pw3\[2\] _01958_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_11600_ channels.pw3\[4\] _03704_ _03705_ _03706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_65_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12580_ _04574_ _04585_ _04586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_65_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_102_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11531_ _03640_ _01880_ _03657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_110_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12636__I _04641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14250_ _06240_ _06248_ _06249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_80_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11462_ channels.accum\[1\]\[16\] _03614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_162_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13201_ _05204_ _05205_ _05206_ _05207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10413_ _02667_ _02668_ _02674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_33_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08759__A2 _01230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14181_ _06070_ _06181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_104_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11393_ channels.accum\[2\]\[11\] _03571_ _03574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13132_ _05135_ _05136_ _05137_ _05138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_10344_ _02603_ _02604_ _02605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_103_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09708__A1 _01807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13063_ net57 _05069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12371__I _04376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10275_ _02535_ _02536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11515__A1 channels.pw1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12014_ channels.env_counter\[1\]\[1\] _04079_ _04081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_109_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16822_ _01766_ _00915_ _00920_ _00919_ _00826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_79_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16753_ _08450_ _00871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_161_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13965_ _05966_ _05963_ _05967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_15704_ channels.exp_periods\[3\]\[4\] _07627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12916_ _04921_ _04917_ _04922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_17_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16684_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[6\] _08244_ _08425_ _08426_
+ _08427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_122_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13896_ _05889_ _05897_ _05898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_122_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16727__B _08459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15635_ _07566_ _07567_ _07568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_150_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12847_ _04476_ _04396_ _04853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_158_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15566_ _07502_ _07503_ _07504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__16509__A2 _08289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12778_ _04783_ _04784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09644__B1 _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17305_ _00375_ clknet_leaf_146_clk channels.accum\[1\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14517_ _06409_ _06489_ _06513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_11729_ channels.atk_dec1\[3\] channels.sus_rel1\[3\] _03785_ _03820_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_127_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15497_ _07439_ _07440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17236_ _00306_ clknet_leaf_170_clk channels.sample1\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14448_ _06435_ _06444_ _06445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_114_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17167_ _00237_ clknet_leaf_146_clk channels.ctrl_reg3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13743__A2 _05746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14379_ _06238_ _06239_ _06377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_168_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09855__I channels.pw2\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16118_ _07991_ _07993_ _07995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_40_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17098_ _00168_ clknet_leaf_98_clk channels.ctrl_reg1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_101_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12281__I _04286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16049_ _07841_ _07754_ _07928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08940_ _01349_ _01405_ _01406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08871_ channels.accum\[0\]\[2\] channels.accum\[1\]\[2\] channels.accum\[2\]\[2\]
+ channels.accum\[3\]\[2\] _01145_ _01159_ _01342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XTAP_TAPCELL_ROW_181_3737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_3748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_232_clk clknet_5_17__leaf_clk clknet_leaf_232_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_159_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09423_ _01814_ _01802_ _01815_ _00139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__14936__I _06909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_179_3699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09354_ _01755_ _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_137_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_47_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10245__A1 _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09285_ channels.lfsr\[1\]\[20\] _01713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11993__A1 _04044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14931__A1 filters.band\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10704__I _02657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10060_ _02334_ _02335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_223_clk clknet_5_20__leaf_clk clknet_leaf_223_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_89_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10720__A2 _02973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15007__I _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13750_ _03269_ _03346_ _05753_ _05754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10962_ _03186_ _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__13670__A1 _04211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12473__A2 _04278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12701_ _04702_ _04704_ _04706_ _04707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_167_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11681__B1 _03771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13681_ _05609_ _05684_ _05614_ _05685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10893_ _03138_ _03141_ _03142_ _00282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15420_ filters.high\[25\] _07369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_127_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12632_ _04613_ _04541_ _04637_ _04594_ _04638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XANTENNA__08844__I _01253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13422__A1 _05405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13422__B2 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12366__I _04371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12563_ _04565_ _04567_ _04569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_15351_ _07295_ _06294_ _07292_ _07306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_80_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12776__A3 _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11514_ _03511_ _03642_ _03646_ _00399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_19_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14302_ _06169_ _06299_ _06300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_80_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12494_ _04288_ _04500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_81_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15282_ filters.high\[13\] _07033_ _06899_ _07243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_108_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16282__B _07740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15714__A3 _03205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09929__A1 _02240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17021_ _00100_ clknet_leaf_231_clk channels.lfsr\[2\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14233_ _06147_ _06156_ _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14922__A1 _05547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11445_ _03602_ _03603_ _01420_ _03604_ _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_145_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14164_ _06082_ _06163_ _06164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_104_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11376_ _03563_ _03557_ _01372_ _03558_ _00344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_104_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15478__A2 _06983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_156_Right_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10614__I _02872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13115_ _05118_ _05119_ _05120_ _05121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_10327_ _01521_ _02381_ _02586_ _02550_ _02587_ _02588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_14095_ _06007_ _06009_ _06094_ _06095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_163_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13046_ _04925_ _05050_ _05051_ _05052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_163_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10258_ _02518_ _02519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_214_clk clknet_5_21__leaf_clk clknet_leaf_214_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_79_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10189_ _01527_ _02448_ _02436_ _02449_ _02450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_16805_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[1\] _00907_ _00909_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17785_ _00855_ clknet_leaf_204_clk channels.exp_periods\[0\]\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14997_ _06959_ _06967_ _06968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_16736_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[5\] _08465_ _08459_ _00860_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_163_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13948_ _05804_ _05948_ _05949_ _05950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_156_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13661__A1 _04562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16457__B _07700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16667_ _08411_ _08412_ _08413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_158_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13879_ _05785_ _05844_ _05881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_88_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15618_ channels.sample2\[8\] _03223_ _07551_ _03232_ _07552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_158_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16598_ _08367_ _08371_ _08372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_56_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10227__A1 _01481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15549_ _07463_ _07488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09093__A1 _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_139_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11180__I _03221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09070_ _01523_ _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_4_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08840__A1 _01308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17219_ _00289_ clknet_leaf_173_clk channels.sample2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_181_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13716__A2 _04753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14913__A1 _06456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11727__A1 channels.sus_rel3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11727__B2 channels.sus_rel2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15469__A2 _07413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09972_ _02101_ _02272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XPHY_EDGE_ROW_123_Right_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10950__A2 _01261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08923_ channels.accum\[0\]\[6\] channels.accum\[1\]\[6\] channels.accum\[2\]\[6\]
+ channels.accum\[3\]\[6\] _01147_ _01162_ _01390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
Xclkbuf_leaf_205_clk clknet_5_23__leaf_clk clknet_leaf_205_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08854_ channels.freq2\[1\] _01274_ _01287_ channels.freq1\[1\] _01326_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_23_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_179_Left_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08785_ _01086_ _01255_ _01258_ channels.ring_outs\[0\] _01259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_46_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13652__A1 _05553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09406_ _01800_ _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_45_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08664__I _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12207__A2 _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10218__A1 channels.pw1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11415__B1 _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09337_ _01739_ _01740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_30_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09268_ _01575_ _01683_ _01698_ _01699_ _00096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_51_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09199_ channels.lfsr\[0\]\[7\] _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11230_ _03439_ _03225_ _03441_ _03442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13183__A3 _05188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11161_ _03376_ _03377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_105_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10112_ channels.ctrl_reg2\[2\] channels.ring_outs\[0\] _01273_ _02373_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11092_ _03283_ _03312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_179_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10043_ _02293_ _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14920_ _06768_ _06884_ _06895_ _06874_ _06886_ _06896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_141_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13891__A1 _04597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12694__A2 _04697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14851_ _06813_ _06824_ _06717_ _06833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13802_ _04728_ _05078_ _05805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17570_ _00640_ clknet_leaf_37_clk filters.low\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13643__A1 _05647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14782_ _06753_ _06757_ _06770_ _06771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11994_ channels.env_counter\[2\]\[12\] _04012_ _04065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16521_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[7\] _08282_ _08252_ _08308_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13733_ _05725_ _05736_ _05737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_82_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10945_ _01320_ _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16452_ _08249_ _08250_ _00733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_27_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13664_ _05582_ _05601_ _05668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10876_ _03117_ _03116_ _03127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15403_ _07350_ _07353_ _07354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12615_ _04618_ _04620_ _04621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16383_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[2\] _08198_ _08199_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13595_ _05591_ _05599_ _05600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_156_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15334_ filters.high\[18\] _06955_ _07290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12546_ _04285_ _04213_ _04305_ _04552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__16345__B1 _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15265_ _01772_ _02056_ _07214_ _07226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12477_ _04404_ _04483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_22_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11709__B2 channels.atk_dec2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17004_ _00083_ clknet_leaf_219_clk channels.lfsr\[2\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_4 _01588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14216_ _06210_ _06214_ _06215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_111_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11428_ _03160_ _01333_ _03594_ _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15196_ _07158_ _07159_ _07160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_123_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14147_ _06143_ _06146_ _06147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_46_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11359_ _03545_ channels.adsr_state\[0\]\[0\] _03552_ _03553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_158_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10932__A2 _02880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15320__A1 _03468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14078_ _05975_ _06078_ _06079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13029_ _05032_ _05034_ _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_20_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08889__A1 _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13882__A1 _04667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10696__A1 _02602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__16820__A1 _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer16 _05287_ net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_179_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer27 net55 net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08570_ _01042_ _01087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xrebuffer38 _07426_ net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_17768_ _00838_ clknet_leaf_203_clk channels.exp_periods\[2\]\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16719_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[6\] _08454_ _08451_ _08455_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17699_ _00769_ clknet_leaf_222_clk channels.lfsr\[0\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_176_3647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_176_3658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09122_ channels.accum\[0\]\[23\] _01560_ _01572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09161__S1 _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09053_ _01507_ _01510_ _01511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__12734__I _04739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14362__A2 _05891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_16__f_clk_I clknet_3_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16639__A1 _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10254__I channels.ch3_env\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10923__A2 _03156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09955_ _02238_ _02257_ _02260_ _00226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_38_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08906_ _01373_ _01371_ _01374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08659__I _01142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09886_ _02179_ _02210_ _02212_ _00205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_148_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12676__A2 _04674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13873__A1 _05846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08837_ _01146_ _01260_ _01309_ _01310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15780__I _07683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16811__A1 _08456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15614__A2 _07543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08768_ _01244_ _00051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_169_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14968__A4 channels.sample2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08699_ _01174_ _01177_ _01182_ _01183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_177_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10730_ _02949_ _02984_ _02985_ _02986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_177_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10661_ _02917_ _02918_ _02919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_94_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09057__A1 _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12400_ _04405_ _04406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_63_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13380_ _04643_ _05054_ _04944_ _05386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_35_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10592_ _02554_ _02601_ _02851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10611__A1 _01705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16878__A1 _00940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12331_ _04335_ _04336_ _04337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_134_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12262_ _04267_ _04268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15050_ _01760_ channels.sample2\[4\] _07019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_181_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_151_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15550__A1 channels.sample3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12364__A1 _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14001_ _05946_ _05955_ _06001_ _06002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_11213_ _03422_ _03224_ _03425_ _03234_ _03426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_31_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12193_ _04198_ _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_102_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10914__A2 _03080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11144_ filters.band\[8\] _03361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_75_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15302__A1 _05968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15952_ _07726_ _07834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11075_ _03281_ _03265_ _03266_ _03296_ _00310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__08569__I _01085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10026_ _02289_ _01943_ _02309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_14903_ _06614_ _06869_ _06860_ _06881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15883_ tt_um_rejunity_sn76489.chan\[1\].attenuation.in _07765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_118_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17622_ _00692_ clknet_leaf_133_clk channels.env_counter\[3\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14834_ _06815_ _06817_ _06818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13616__A1 _03383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17553_ _00623_ clknet_leaf_25_clk filters.low\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_158_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14765_ _03472_ _06755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_11977_ _04019_ _04050_ _04051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_158_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16504_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[4\] _08289_ _08291_ _08293_
+ _08294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_13716_ _04802_ _04753_ _05720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17484_ _00554_ clknet_leaf_244_clk filters.band\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10928_ _01460_ _03164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14696_ _03412_ _03378_ _06690_ _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_50_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16435_ _08235_ _08236_ _08237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09048__A1 channels.freq2\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10339__I _02569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13647_ _05547_ _05651_ _05652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09048__B2 channels.freq1\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10859_ _03089_ _03090_ _03111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_116_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09599__A2 net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16366_ _03964_ _08184_ _08186_ _00711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_171_3555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13578_ _05467_ _05317_ _05473_ _05583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_171_3566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16869__A1 _00940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15317_ _07260_ _07262_ _07275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12529_ _04333_ _04535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16297_ channels.env_counter\[3\]\[4\] _08146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_140_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_132_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_132_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15248_ _07207_ _07208_ _07209_ _07210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_10_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15179_ _03373_ _07064_ _07143_ _07089_ _00567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_22_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16897__S _00975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15844__A2 _07721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09740_ _01756_ _02110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08479__I _01008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
.ends

