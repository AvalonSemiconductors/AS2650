// This is the unpowered netlist.
module timers (bus_cyc,
    bus_we,
    irq1,
    irq2,
    irq5,
    pwm0,
    pwm1,
    pwm2,
    rst,
    tmr0_clk,
    tmr0_o,
    tmr1_clk,
    tmr1_o,
    wb_clk_i,
    addr,
    data_in,
    data_out);
 input bus_cyc;
 input bus_we;
 output irq1;
 output irq2;
 output irq5;
 output pwm0;
 output pwm1;
 output pwm2;
 input rst;
 input tmr0_clk;
 output tmr0_o;
 input tmr1_clk;
 output tmr1_o;
 input wb_clk_i;
 input [5:0] addr;
 input [7:0] data_in;
 output [7:0] data_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0__leaf_wb_clk_i;
 wire clknet_3_1__leaf_wb_clk_i;
 wire clknet_3_2__leaf_wb_clk_i;
 wire clknet_3_3__leaf_wb_clk_i;
 wire clknet_3_4__leaf_wb_clk_i;
 wire clknet_3_5__leaf_wb_clk_i;
 wire clknet_3_6__leaf_wb_clk_i;
 wire clknet_3_7__leaf_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_57_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_60_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_62_wb_clk_i;
 wire clknet_leaf_63_wb_clk_i;
 wire clknet_leaf_64_wb_clk_i;
 wire clknet_leaf_66_wb_clk_i;
 wire clknet_leaf_67_wb_clk_i;
 wire clknet_leaf_69_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_70_wb_clk_i;
 wire clknet_leaf_71_wb_clk_i;
 wire clknet_leaf_72_wb_clk_i;
 wire clknet_leaf_73_wb_clk_i;
 wire clknet_leaf_74_wb_clk_i;
 wire clknet_leaf_76_wb_clk_i;
 wire clknet_leaf_77_wb_clk_i;
 wire clknet_leaf_78_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_81_wb_clk_i;
 wire clknet_leaf_82_wb_clk_i;
 wire clknet_leaf_83_wb_clk_i;
 wire clknet_leaf_84_wb_clk_i;
 wire clknet_leaf_85_wb_clk_i;
 wire clknet_leaf_86_wb_clk_i;
 wire clknet_leaf_87_wb_clk_i;
 wire clknet_leaf_88_wb_clk_i;
 wire clknet_leaf_89_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_90_wb_clk_i;
 wire clknet_leaf_91_wb_clk_i;
 wire clknet_leaf_92_wb_clk_i;
 wire clknet_leaf_93_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire last_tmr0_clk;
 wire last_tmr1_clk;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire \pw0[0] ;
 wire \pw0[1] ;
 wire \pw0[2] ;
 wire \pw0[3] ;
 wire \pw0[4] ;
 wire \pw0[5] ;
 wire \pw0[6] ;
 wire \pw0[7] ;
 wire \pw1[0] ;
 wire \pw1[1] ;
 wire \pw1[2] ;
 wire \pw1[3] ;
 wire \pw1[4] ;
 wire \pw1[5] ;
 wire \pw1[6] ;
 wire \pw1[7] ;
 wire \pw2[0] ;
 wire \pw2[1] ;
 wire \pw2[2] ;
 wire \pw2[3] ;
 wire \pw2[4] ;
 wire \pw2[5] ;
 wire \pw2[6] ;
 wire \pw2[7] ;
 wire \pwm_ctr0[0] ;
 wire \pwm_ctr0[1] ;
 wire \pwm_ctr0[2] ;
 wire \pwm_ctr0[3] ;
 wire \pwm_ctr0[4] ;
 wire \pwm_ctr0[5] ;
 wire \pwm_ctr0[6] ;
 wire \pwm_ctr0[7] ;
 wire \pwm_ctr1[0] ;
 wire \pwm_ctr1[1] ;
 wire \pwm_ctr1[2] ;
 wire \pwm_ctr1[3] ;
 wire \pwm_ctr1[4] ;
 wire \pwm_ctr1[5] ;
 wire \pwm_ctr1[6] ;
 wire \pwm_ctr1[7] ;
 wire \pwm_ctr2[0] ;
 wire \pwm_ctr2[1] ;
 wire \pwm_ctr2[2] ;
 wire \pwm_ctr2[3] ;
 wire \pwm_ctr2[4] ;
 wire \pwm_ctr2[5] ;
 wire \pwm_ctr2[6] ;
 wire \pwm_ctr2[7] ;
 wire \settings[0] ;
 wire \settings[1] ;
 wire \settings[2] ;
 wire \t0_capture[0] ;
 wire \t0_capture[10] ;
 wire \t0_capture[11] ;
 wire \t0_capture[12] ;
 wire \t0_capture[13] ;
 wire \t0_capture[14] ;
 wire \t0_capture[15] ;
 wire \t0_capture[1] ;
 wire \t0_capture[2] ;
 wire \t0_capture[3] ;
 wire \t0_capture[4] ;
 wire \t0_capture[5] ;
 wire \t0_capture[6] ;
 wire \t0_capture[7] ;
 wire \t0_capture[8] ;
 wire \t0_capture[9] ;
 wire \t0_top[0] ;
 wire \t0_top[10] ;
 wire \t0_top[11] ;
 wire \t0_top[12] ;
 wire \t0_top[13] ;
 wire \t0_top[14] ;
 wire \t0_top[15] ;
 wire \t0_top[1] ;
 wire \t0_top[2] ;
 wire \t0_top[3] ;
 wire \t0_top[4] ;
 wire \t0_top[5] ;
 wire \t0_top[6] ;
 wire \t0_top[7] ;
 wire \t0_top[8] ;
 wire \t0_top[9] ;
 wire \t0pre[0] ;
 wire \t0pre[10] ;
 wire \t0pre[11] ;
 wire \t0pre[12] ;
 wire \t0pre[13] ;
 wire \t0pre[14] ;
 wire \t0pre[15] ;
 wire \t0pre[1] ;
 wire \t0pre[2] ;
 wire \t0pre[3] ;
 wire \t0pre[4] ;
 wire \t0pre[5] ;
 wire \t0pre[6] ;
 wire \t0pre[7] ;
 wire \t0pre[8] ;
 wire \t0pre[9] ;
 wire \t0pre_counter[0] ;
 wire \t0pre_counter[10] ;
 wire \t0pre_counter[11] ;
 wire \t0pre_counter[12] ;
 wire \t0pre_counter[13] ;
 wire \t0pre_counter[14] ;
 wire \t0pre_counter[15] ;
 wire \t0pre_counter[1] ;
 wire \t0pre_counter[2] ;
 wire \t0pre_counter[3] ;
 wire \t0pre_counter[4] ;
 wire \t0pre_counter[5] ;
 wire \t0pre_counter[6] ;
 wire \t0pre_counter[7] ;
 wire \t0pre_counter[8] ;
 wire \t0pre_counter[9] ;
 wire \t1_capture[0] ;
 wire \t1_capture[10] ;
 wire \t1_capture[11] ;
 wire \t1_capture[12] ;
 wire \t1_capture[13] ;
 wire \t1_capture[14] ;
 wire \t1_capture[15] ;
 wire \t1_capture[1] ;
 wire \t1_capture[2] ;
 wire \t1_capture[3] ;
 wire \t1_capture[4] ;
 wire \t1_capture[5] ;
 wire \t1_capture[6] ;
 wire \t1_capture[7] ;
 wire \t1_capture[8] ;
 wire \t1_capture[9] ;
 wire \t1_top[0] ;
 wire \t1_top[10] ;
 wire \t1_top[11] ;
 wire \t1_top[12] ;
 wire \t1_top[13] ;
 wire \t1_top[14] ;
 wire \t1_top[15] ;
 wire \t1_top[1] ;
 wire \t1_top[2] ;
 wire \t1_top[3] ;
 wire \t1_top[4] ;
 wire \t1_top[5] ;
 wire \t1_top[6] ;
 wire \t1_top[7] ;
 wire \t1_top[8] ;
 wire \t1_top[9] ;
 wire \t1pre[0] ;
 wire \t1pre[10] ;
 wire \t1pre[11] ;
 wire \t1pre[12] ;
 wire \t1pre[13] ;
 wire \t1pre[14] ;
 wire \t1pre[15] ;
 wire \t1pre[1] ;
 wire \t1pre[2] ;
 wire \t1pre[3] ;
 wire \t1pre[4] ;
 wire \t1pre[5] ;
 wire \t1pre[6] ;
 wire \t1pre[7] ;
 wire \t1pre[8] ;
 wire \t1pre[9] ;
 wire \t1pre_counter[0] ;
 wire \t1pre_counter[10] ;
 wire \t1pre_counter[11] ;
 wire \t1pre_counter[12] ;
 wire \t1pre_counter[13] ;
 wire \t1pre_counter[14] ;
 wire \t1pre_counter[15] ;
 wire \t1pre_counter[1] ;
 wire \t1pre_counter[2] ;
 wire \t1pre_counter[3] ;
 wire \t1pre_counter[4] ;
 wire \t1pre_counter[5] ;
 wire \t1pre_counter[6] ;
 wire \t1pre_counter[7] ;
 wire \t1pre_counter[8] ;
 wire \t1pre_counter[9] ;
 wire \t2_capture[0] ;
 wire \t2_capture[10] ;
 wire \t2_capture[11] ;
 wire \t2_capture[12] ;
 wire \t2_capture[13] ;
 wire \t2_capture[14] ;
 wire \t2_capture[15] ;
 wire \t2_capture[1] ;
 wire \t2_capture[2] ;
 wire \t2_capture[3] ;
 wire \t2_capture[4] ;
 wire \t2_capture[5] ;
 wire \t2_capture[6] ;
 wire \t2_capture[7] ;
 wire \t2_capture[8] ;
 wire \t2_capture[9] ;
 wire \t2_top[0] ;
 wire \t2_top[10] ;
 wire \t2_top[11] ;
 wire \t2_top[12] ;
 wire \t2_top[13] ;
 wire \t2_top[14] ;
 wire \t2_top[15] ;
 wire \t2_top[1] ;
 wire \t2_top[2] ;
 wire \t2_top[3] ;
 wire \t2_top[4] ;
 wire \t2_top[5] ;
 wire \t2_top[6] ;
 wire \t2_top[7] ;
 wire \t2_top[8] ;
 wire \t2_top[9] ;
 wire \t2pre[0] ;
 wire \t2pre[10] ;
 wire \t2pre[11] ;
 wire \t2pre[12] ;
 wire \t2pre[13] ;
 wire \t2pre[14] ;
 wire \t2pre[15] ;
 wire \t2pre[1] ;
 wire \t2pre[2] ;
 wire \t2pre[3] ;
 wire \t2pre[4] ;
 wire \t2pre[5] ;
 wire \t2pre[6] ;
 wire \t2pre[7] ;
 wire \t2pre[8] ;
 wire \t2pre[9] ;
 wire \t2pre_counter[0] ;
 wire \t2pre_counter[10] ;
 wire \t2pre_counter[11] ;
 wire \t2pre_counter[12] ;
 wire \t2pre_counter[13] ;
 wire \t2pre_counter[14] ;
 wire \t2pre_counter[15] ;
 wire \t2pre_counter[1] ;
 wire \t2pre_counter[2] ;
 wire \t2pre_counter[3] ;
 wire \t2pre_counter[4] ;
 wire \t2pre_counter[5] ;
 wire \t2pre_counter[6] ;
 wire \t2pre_counter[7] ;
 wire \t2pre_counter[8] ;
 wire \t2pre_counter[9] ;
 wire \temp[0] ;
 wire \temp[1] ;
 wire \temp[2] ;
 wire \temp[3] ;
 wire \temp[4] ;
 wire \temp[5] ;
 wire \temp[6] ;
 wire \temp[7] ;
 wire \timer0[0] ;
 wire \timer0[10] ;
 wire \timer0[11] ;
 wire \timer0[12] ;
 wire \timer0[13] ;
 wire \timer0[14] ;
 wire \timer0[15] ;
 wire \timer0[1] ;
 wire \timer0[2] ;
 wire \timer0[3] ;
 wire \timer0[4] ;
 wire \timer0[5] ;
 wire \timer0[6] ;
 wire \timer0[7] ;
 wire \timer0[8] ;
 wire \timer0[9] ;
 wire \timer1[0] ;
 wire \timer1[10] ;
 wire \timer1[11] ;
 wire \timer1[12] ;
 wire \timer1[13] ;
 wire \timer1[14] ;
 wire \timer1[15] ;
 wire \timer1[1] ;
 wire \timer1[2] ;
 wire \timer1[3] ;
 wire \timer1[4] ;
 wire \timer1[5] ;
 wire \timer1[6] ;
 wire \timer1[7] ;
 wire \timer1[8] ;
 wire \timer1[9] ;
 wire \timer2[0] ;
 wire \timer2[10] ;
 wire \timer2[11] ;
 wire \timer2[12] ;
 wire \timer2[13] ;
 wire \timer2[14] ;
 wire \timer2[15] ;
 wire \timer2[1] ;
 wire \timer2[2] ;
 wire \timer2[3] ;
 wire \timer2[4] ;
 wire \timer2[5] ;
 wire \timer2[6] ;
 wire \timer2[7] ;
 wire \timer2[8] ;
 wire \timer2[9] ;
 wire tmr0_ext;
 wire tmr1_ext;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2105__A1 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2107__A1 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2109__A1 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2110__I (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2111__C (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2112__A1 (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__I (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2115__I (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2117__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__C (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2120__A1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2121__C (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2123__C (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2125__I (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2128__A1 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2131__A1 (.I(\temp[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2133__A1 (.I(\temp[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2135__A1 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2136__I (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2139__A1 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2142__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2144__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2146__A1 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2147__I (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2149__A1 (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2149__A2 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2150__A1 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2150__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2151__A1 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2152__A1 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2153__A1 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2153__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2154__A1 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2154__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2155__A1 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__A1 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2159__A1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2159__A2 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2160__I (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2161__I (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__I (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__I (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2176__A1 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2176__A3 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2178__A3 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2179__A2 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2180__A2 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2181__A2 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2183__A1 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2188__B (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2197__A1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2199__A1 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2201__A2 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__A1 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2207__B (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2211__A1 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2213__A1 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2216__A1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__A1 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2220__A2 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__A1 (.I(\pw0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2222__A1 (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2222__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2224__A1 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2225__B (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2228__I (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2229__A1 (.I(\pw0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2230__A1 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2232__A1 (.I(\pw0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2233__A1 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2234__A1 (.I(\pw0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__A1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__B (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__A1 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__C (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2240__A1 (.I(\pw0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2241__A1 (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2242__A1 (.I(\pw0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2243__A1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2244__A1 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2245__A1 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2245__C (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2246__A2 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2247__A1 (.I(\pw1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2249__I (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2250__A1 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2250__A2 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2251__B (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2252__I (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__I (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2254__I (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2255__A1 (.I(\pw1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2256__A1 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__A1 (.I(\pw1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2258__A1 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2259__A1 (.I(\pw1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2260__A1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2260__A2 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2261__B (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2263__I (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2265__A1 (.I(\pw1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2266__A1 (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2267__A1 (.I(\pw1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2268__A1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2269__A1 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2269__A2 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2270__A2 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2270__C (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2271__A2 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2273__A1 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2274__A1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2276__I (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2277__I (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2278__I (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2279__A1 (.I(\pw2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__A1 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__A1 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2283__A1 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2286__A1 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2287__A1 (.I(\pw2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2287__A2 (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2288__A1 (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2289__A1 (.I(\pw2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2289__A2 (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__A1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2291__A1 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2292__A1 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2292__C (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2295__A1 (.I(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2296__I (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2297__A1 (.I(\temp[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2300__A1 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2300__A2 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__B (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2302__I (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2303__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2304__I (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2305__A1 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2306__A2 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2306__B (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2307__A1 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2307__A2 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__I (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2310__A1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2311__A1 (.I(\temp[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2312__A1 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2312__A2 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2313__B (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2315__A1 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2316__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2317__A1 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2318__A1 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2319__A1 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2319__C (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2321__I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__I (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2323__I (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2324__I (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2325__A2 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2328__I (.I(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2331__A1 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__I (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2336__A1 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2339__A1 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__A1 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__A1 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2349__A1 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2351__I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2353__I (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2355__B (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2359__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2361__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2362__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2363__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2364__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2369__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2370__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2373__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__A2 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__B2 (.I(\t0pre[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2384__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__A1 (.I(\t0pre[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__B1 (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__B2 (.I(\settings[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2393__I (.I(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2399__A1 (.I(\t1_capture[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2399__A2 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2399__B1 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2399__B2 (.I(\t2_top[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2402__I (.I(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__A1 (.I(\t2pre[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__A2 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__B2 (.I(\t2_capture[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2412__I (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__A1 (.I(\t0_top[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2414__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2414__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2415__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__B (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__A2 (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__I (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2426__A1 (.I(\t1pre[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2426__B1 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2426__B2 (.I(\t0_capture[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2426__C1 (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2426__C2 (.I(\t2_top[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2431__I (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2432__A1 (.I(\pw0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2432__A2 (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__A4 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__A1 (.I(\t0_top[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__B2 (.I(\t1_top[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2444__I (.I(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2446__B2 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2451__A2 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2451__B2 (.I(\t2pre[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__I (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2456__A1 (.I(\t1_top[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2456__B2 (.I(\pw1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2457__A2 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2460__B2 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2463__I (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__A1 (.I(\t1_top[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__B2 (.I(\t2pre[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__A1 (.I(\t0_top[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2471__A1 (.I(\t1_capture[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2472__I (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2473__I (.I(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2475__A1 (.I(\pw0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2475__B2 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__A2 (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2477__I (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__I (.I(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__A1 (.I(\pw2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2482__I (.I(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__B2 (.I(\t1pre[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__A1 (.I(\t2_top[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__A2 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__B2 (.I(\t0_capture[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__C1 (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A2 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__A1 (.I(\t0_top[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__B1 (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__B2 (.I(\t2_top[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__A1 (.I(\t0pre[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2490__A1 (.I(\pw1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2490__B2 (.I(\t1_top[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2491__A1 (.I(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2491__A3 (.I(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2492__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__A1 (.I(\t1_top[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__B2 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2496__A1 (.I(\t0_top[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2496__B2 (.I(\t2_capture[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__A1 (.I(\t1_capture[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__B2 (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A1 (.I(\pw0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__B2 (.I(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__A2 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__A1 (.I(\t1pre[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__B2 (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__A1 (.I(\t2_top[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__A2 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__B2 (.I(\t0_capture[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__C1 (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__I (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__I (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2510__B2 (.I(\t2_top[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__A1 (.I(\t0pre[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__A3 (.I(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2515__A1 (.I(\pw1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2515__B2 (.I(\t1_top[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__A1 (.I(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__A3 (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__A1 (.I(\t1_top[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__B2 (.I(\t2pre[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__A1 (.I(\t0_top[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__B2 (.I(\t2_capture[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__A1 (.I(\t1_capture[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__B2 (.I(\t0pre[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2522__A1 (.I(\pw0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2522__B2 (.I(\t2pre[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__A2 (.I(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2526__B2 (.I(\t1pre[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2527__A1 (.I(\t2_top[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2527__A2 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2527__B2 (.I(\t0_capture[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2527__C1 (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2527__C2 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__B2 (.I(\t2_top[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2532__A1 (.I(\t0pre[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__A3 (.I(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2534__A1 (.I(\pw1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2534__B2 (.I(\t1_top[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2535__A1 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2535__A3 (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A1 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__A1 (.I(\t1_top[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__B2 (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2540__A1 (.I(\t0_top[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2540__B2 (.I(\t2_capture[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2542__A1 (.I(\t1_capture[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2542__B2 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2543__I (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2545__A2 (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__B2 (.I(\t1pre[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2549__A1 (.I(\t2_top[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2549__B2 (.I(\t0_capture[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2549__C2 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2553__B2 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2554__A1 (.I(\t0pre[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2555__A3 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2555__A4 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2556__A1 (.I(\pw1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2556__B2 (.I(\t1_top[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__A2 (.I(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__A3 (.I(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2558__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2560__A1 (.I(\t1_top[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2560__B2 (.I(\t2pre[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2561__A1 (.I(\t0_top[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2561__B2 (.I(\t2_capture[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2563__A2 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2563__B2 (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__A1 (.I(\pw0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__B1 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__A2 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2566__A1 (.I(\pw2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2566__B1 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2568__B2 (.I(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2569__A1 (.I(\t2_top[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2569__B1 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2569__B2 (.I(\t0_capture[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2569__C2 (.I(tmr0_ext));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__B2 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2573__A1 (.I(\t0pre[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2574__A3 (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2574__A4 (.I(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__A1 (.I(\pw1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__B2 (.I(\t1_top[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__A1 (.I(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__A2 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__A3 (.I(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2577__A1 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2580__A1 (.I(\t1_top[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2580__B2 (.I(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2581__A1 (.I(\t0_top[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2581__B2 (.I(\t2_capture[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__A1 (.I(\t1_capture[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__A2 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__B2 (.I(\t0pre[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__A1 (.I(\pw0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__B1 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2584__A2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2585__A1 (.I(\pw2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2585__B1 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2587__B2 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__A1 (.I(\t2_top[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__B1 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__B2 (.I(\t0_capture[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__A2 (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__B1 (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2591__A1 (.I(\t0pre[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2592__A3 (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__A1 (.I(\pw1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__B2 (.I(\t1_top[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__A1 (.I(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__A2 (.I(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__A3 (.I(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2595__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2598__A1 (.I(\t0_top[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2598__B2 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__A1 (.I(\t2pre[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__A2 (.I(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__B1 (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__B2 (.I(\t2_top[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2600__B1 (.I(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2600__B2 (.I(\t1_capture[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2602__A1 (.I(\t0pre[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2602__B2 (.I(\t2_capture[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__A2 (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__B1 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2604__A1 (.I(\t2_top[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2604__B1 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2604__B2 (.I(\t0_capture[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2605__A1 (.I(\t1_top[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2605__A2 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2605__B2 (.I(\t2_capture[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2606__A1 (.I(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2606__A2 (.I(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2607__A1 (.I(\t0_top[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2607__B2 (.I(\t0pre[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__A1 (.I(\t1_top[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__A1 (.I(\pw1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__B1 (.I(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__B2 (.I(\t1pre[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__A1 (.I(\pw0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__B1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2613__A1 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__I (.I(\settings[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2616__I (.I(\t0pre[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2625__A2 (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__I (.I(\t0pre[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__A2 (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2643__I (.I(\t0pre[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2646__A1 (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__A2 (.I(\t0pre[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__A1 (.I(\t0pre[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__A1 (.I(\t0pre[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2650__I (.I(\t0pre[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2654__I (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2660__A1 (.I(\t0pre[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2664__A1 (.I(\t0pre[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2664__B2 (.I(\t0pre[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2665__I (.I(\t0pre[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__I (.I(\t0pre[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__B (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__A1 (.I(\t0pre[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__B2 (.I(\t0pre[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2675__I (.I(\t0pre[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2688__A1 (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2688__B2 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2691__A1 (.I(\t0pre[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2691__B2 (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__I (.I(\t0pre[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2699__A1 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2709__A1 (.I(\t0pre[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2709__B2 (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2713__A2 (.I(\t0pre[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2715__A1 (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2716__A1 (.I(\t0pre[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2721__A1 (.I(\t0pre[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__I (.I(\t0pre[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2727__A1 (.I(\t0pre[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__A2 (.I(\t0pre[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__I (.I(tmr0_ext));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2739__I (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__I (.I(\t0_top[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__I (.I(\t0_top[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__I (.I(\timer0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2746__I (.I(\t0_top[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2747__I (.I(\t0_top[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2748__I (.I(\timer0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2750__I (.I(\t0_top[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2753__A1 (.I(\t0_top[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2753__B (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2753__C (.I(\t0_top[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2754__I (.I(\timer0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2755__A1 (.I(\t0_top[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2755__B2 (.I(\t0_top[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2756__A1 (.I(\t0_top[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2756__A2 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2757__A2 (.I(\timer0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2758__A1 (.I(\t0_top[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2758__B1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2758__B2 (.I(\t0_top[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2759__A2 (.I(\timer0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2759__B1 (.I(\timer0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__A1 (.I(\t0_top[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__A2 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__B1 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__B2 (.I(\t0_top[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2761__A2 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2761__B1 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2765__B1 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2767__I (.I(\timer0[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2768__A1 (.I(\t0_top[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2768__A2 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2768__B1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2768__B2 (.I(\t0_top[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2771__A2 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2771__B1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2771__B2 (.I(\t0_top[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2773__I (.I(\t0_top[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2775__A2 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2776__A2 (.I(\timer0[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2777__I (.I(\timer0[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2778__A1 (.I(\t0_top[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2778__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2780__A2 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2781__I (.I(\t0_top[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__A2 (.I(\timer0[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2785__I (.I(\timer0[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2786__A2 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2786__B1 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2788__A2 (.I(\timer0[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__A2 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2800__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2808__I (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2809__A1 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2809__A2 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2809__C (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2810__A2 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2811__I (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2813__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2814__A1 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2814__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2817__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2817__B (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2824__A2 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__A2 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2837__A1 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2847__A1 (.I(\t1pre[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2855__A1 (.I(\t1pre[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2861__I (.I(\t1pre[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2864__B2 (.I(\t1pre[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2872__A1 (.I(\t1pre[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2875__A2 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2876__A1 (.I(\t1pre[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2877__A1 (.I(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2880__A1 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2880__B2 (.I(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2881__A1 (.I(\t1pre[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2881__B2 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2888__A1 (.I(\t1pre[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__A1 (.I(\t1pre[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__B2 (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2899__A1 (.I(\t1pre[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2902__A1 (.I(\t1pre[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2904__A1 (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2905__A1 (.I(\t1pre[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2915__B2 (.I(\t1pre[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2922__A2 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2923__A2 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2929__I (.I(\timer1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__A1 (.I(\t1_top[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__A2 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2931__I (.I(\t1_top[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2934__A1 (.I(\t1_top[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2935__I (.I(\t1_top[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2937__I (.I(\t1_top[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2942__A1 (.I(\t1_top[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2942__B2 (.I(\t1_top[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2945__A1 (.I(\t1_top[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2945__B2 (.I(\t1_top[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2947__A1 (.I(\t1_top[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2947__B2 (.I(\t1_top[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2949__I (.I(\t1_top[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2953__I (.I(\t1_top[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2954__A2 (.I(\timer1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2957__I (.I(\t1_top[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2960__I (.I(\t1_top[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2962__I (.I(\t1_top[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2963__A2 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2963__B (.I(\timer1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2964__A1 (.I(\t1_top[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2964__A2 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2964__B1 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2964__B2 (.I(\t1_top[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2966__A1 (.I(\t1_top[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2966__A2 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2966__B1 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2966__B2 (.I(\t1_top[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2967__A1 (.I(\t1_top[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2967__A2 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2969__I (.I(\t1_top[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2971__B1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2973__A1 (.I(\t1_top[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2973__A2 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2973__C1 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2973__C2 (.I(\t1_top[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2976__A1 (.I(\t1_top[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2976__A2 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2976__B1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2976__B2 (.I(\t1_top[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2980__A1 (.I(\t1_top[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2980__B2 (.I(\t1_top[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2980__C2 (.I(\t1_top[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2986__A1 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2986__A2 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2987__I1 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2987__S (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2988__A1 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2990__A2 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2990__B (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2991__A2 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2993__A2 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2994__A1 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2997__A1 (.I(\pw0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2997__B (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3000__I (.I(\pw0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3002__A1 (.I(\pw0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3003__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3007__A1 (.I(\pw0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3007__B2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3007__C1 (.I(\pw0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3008__I (.I(\pw0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3009__I (.I(\pw0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3010__B2 (.I(\pw0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3011__A1 (.I(\pw0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3011__B2 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3012__A1 (.I(\pw0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3019__A1 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3019__B (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3022__A1 (.I(\pw1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3023__I (.I(\pw1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3025__I (.I(\pw1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3027__A1 (.I(\pw1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3032__A1 (.I(\pw1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3032__C1 (.I(\pw1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3033__I (.I(\pw1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3034__I (.I(\pw1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3035__B2 (.I(\pw1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3036__A1 (.I(\pw1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3037__A1 (.I(\pw1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3044__A1 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3044__B (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3047__I (.I(\pw2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3048__A1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3048__B2 (.I(\pw2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3052__A1 (.I(\pw2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3052__B2 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3054__A1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3057__B2 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3061__A1 (.I(\pw2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3061__B (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__B2 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__C1 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3063__A1 (.I(\pw2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3064__A2 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3067__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3070__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3071__A2 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3071__A3 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3072__A1 (.I(\settings[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3073__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3074__I (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3075__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3075__A2 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3075__A3 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3077__A1 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3078__B (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3079__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3081__B (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3082__A1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3083__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3086__B (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3087__A1 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3088__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3090__A1 (.I(tmr0_ext));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3090__B (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3091__A1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3092__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3093__A1 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3095__A1 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3095__C (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3104__I (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3118__B2 (.I(\t2pre[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3122__I (.I(\t2pre[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3128__A2 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3145__A1 (.I(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3145__B2 (.I(\t2pre[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3146__I (.I(\t2pre[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3149__B2 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3154__I (.I(\t2pre[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3155__B2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3157__A1 (.I(\t2pre[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3164__I (.I(\t2pre[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3182__A1 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3182__C2 (.I(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3188__B2 (.I(\t2pre[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3190__A1 (.I(\t2pre[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3191__A1 (.I(\t2pre[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3191__B2 (.I(\t2pre[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3193__A1 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3195__A1 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3195__B2 (.I(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3197__A1 (.I(\t2pre[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3197__B2 (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3198__A1 (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3198__B2 (.I(\t2pre[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3202__A1 (.I(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3202__B2 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3212__A1 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3213__A1 (.I(\t2pre[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__I (.I(\t2_top[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3222__A2 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3226__B1 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3226__B2 (.I(\t2_top[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3227__I (.I(\t2_top[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3230__I (.I(\t2_top[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3232__I (.I(\t2_top[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__I (.I(\t2_top[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3239__A1 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3239__A2 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3239__B1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3239__B2 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3246__I (.I(\t2_top[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3249__I (.I(\t2_top[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3252__I (.I(\t2_top[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3254__I (.I(\t2_top[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3255__A2 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3255__B1 (.I(\timer2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3256__I (.I(\t2_top[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3258__I (.I(\t2_top[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3262__I (.I(\t2_top[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3265__I (.I(\t2_top[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3267__A1 (.I(\t2_top[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3269__A1 (.I(\t2_top[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3270__I (.I(\timer2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3272__A1 (.I(\t2_top[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3272__A2 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3272__B2 (.I(\t2_top[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3275__A1 (.I(\t2_top[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3275__A2 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3277__A1 (.I(\t2_top[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3277__A2 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3281__A1 (.I(\t2_top[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3281__A2 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3283__A1 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3283__A2 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3283__B1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3283__B2 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3286__A1 (.I(\t2_top[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3286__B1 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3286__B2 (.I(\t2_top[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3297__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3297__A2 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__B1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__C (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3301__A2 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3301__B (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3303__A1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3305__A1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3305__A2 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3309__A3 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3310__I (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3313__I (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3314__I (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3315__A1 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3317__I (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3319__A1 (.I(\temp[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3320__A1 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3323__A1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3323__A2 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3324__I (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3326__I (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3329__I (.I(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3331__A1 (.I(\timer0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3333__I (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3334__A1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3334__A2 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3335__A1 (.I(\timer0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3335__C (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3338__A1 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3341__I (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3343__C (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3344__I (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3345__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3348__I (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3349__I (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3350__A1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3350__C (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3351__I (.I(\temp[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3352__A1 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3352__A2 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3353__I (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3355__I (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3356__A1 (.I(\timer0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3358__A1 (.I(\timer0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3358__C (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3360__I (.I(\temp[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3361__A1 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3362__A1 (.I(\timer0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3363__A1 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3363__C (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3364__I (.I(\temp[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3366__A1 (.I(\timer0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3367__A1 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3368__B (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3369__A1 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3370__I (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3371__I (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3372__A1 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3374__A1 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3375__A1 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3376__A1 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3377__B (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3380__A1 (.I(\timer0[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3380__A3 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__A1 (.I(\timer0[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__C (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3383__A1 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3383__A2 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3384__I (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3385__I (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3386__B (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3388__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3390__A1 (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3393__A1 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3393__A2 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3395__A1 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3396__A1 (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3398__A1 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3400__A1 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3401__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3402__B (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3404__B (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3405__A1 (.I(\timer0[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3405__A2 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3405__A3 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3407__A1 (.I(\timer0[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3407__C (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3408__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3410__A1 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3410__A2 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3411__B (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3413__A1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3414__B2 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3416__I (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3417__A1 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3417__C (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3423__A1 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3424__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3424__C (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3425__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3426__A1 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3427__A2 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3428__A1 (.I(\timer0[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3429__B (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__I (.I(\temp[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__A3 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__I (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3434__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3435__I (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3437__A1 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3437__A2 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3438__I (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3439__I (.I(\timer1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3440__B (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3441__A2 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3443__I (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3445__A1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3446__I (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3447__A1 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3447__A3 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3448__I (.I(\timer1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__I (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3450__I (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3451__I (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3453__A1 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3453__A2 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3453__A3 (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3453__B (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3456__I (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3457__A1 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3460__A2 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3462__A1 (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__I (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3467__A1 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3469__I (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__A1 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3478__A1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3480__A1 (.I(\temp[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3481__A1 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3481__A2 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3481__A3 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3483__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3485__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3491__I (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3492__A1 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3493__A1 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3499__A1 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3500__A1 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3501__A1 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__A3 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3505__A1 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3505__B (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3507__I (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3509__I (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3511__A1 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3511__A3 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3514__C (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3515__A1 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3520__A1 (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3526__A1 (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3527__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__A1 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__A3 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3539__A1 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__A1 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__C (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3549__I (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3550__C (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3551__A1 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3553__A1 (.I(\timer1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3553__C (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3554__I (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3555__B (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__I (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__I (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3561__I (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3562__A1 (.I(\t0_capture[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3562__B (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3563__A1 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__A1 (.I(\t0_capture[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__B (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__A1 (.I(\t0_capture[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__A1 (.I(\t0_capture[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3570__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3571__I (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3572__I (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3573__A1 (.I(\t0_capture[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3575__A1 (.I(\t0_capture[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3576__A1 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3577__I (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3579__A1 (.I(\t0_capture[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3579__B (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3580__A1 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__I (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3582__A1 (.I(\t0_capture[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3582__B (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3584__I (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3586__I (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3588__B (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__A1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3590__B (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3591__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3594__A1 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3595__A3 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__A2 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__I (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__B (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3602__A1 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3606__A1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3608__A1 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3611__A1 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3613__A1 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__A1 (.I(\t1_capture[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3617__A1 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__A1 (.I(\t1_capture[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__A1 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__A1 (.I(\t1_capture[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__A1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3623__A1 (.I(\t1_capture[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3623__A2 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3624__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3624__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__B (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__A1 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__A1 (.I(\t1_capture[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__A1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3633__A1 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__I (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__I (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__A1 (.I(\t1_capture[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3640__I (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__I (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3643__I (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3648__A2 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3649__I (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3650__A2 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__B (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3652__I (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__B (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3655__B (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3657__I (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3658__I (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__A1 (.I(\t1_capture[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__B (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__A1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__A1 (.I(\t2_capture[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__B (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3665__A2 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3667__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3667__A2 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__B (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__I (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__A1 (.I(\t2_capture[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__A1 (.I(\t2_capture[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__I (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3677__I (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__A1 (.I(\t2_capture[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3679__A1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__A1 (.I(\t2_capture[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__A1 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3682__I (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3683__A1 (.I(\t2_capture[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__A1 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3685__A1 (.I(\t2_capture[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3686__A1 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__I (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3688__I (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3690__A1 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__A1 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__A2 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__B (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3697__A1 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3697__A2 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3698__B (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__A1 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3702__I (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3704__A1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3706__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3707__A2 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3708__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3708__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3709__A1 (.I(\t2_capture[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3709__A2 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3710__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3712__A2 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3714__A1 (.I(\t0pre[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3715__I (.I(\temp[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3720__A1 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3721__B (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__I (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3727__I (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__A1 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3731__A1 (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3733__I (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3735__A1 (.I(\t0pre[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3736__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__A1 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3738__I (.I(\temp[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3739__A1 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3742__I (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__A1 (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__A1 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__I (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__A1 (.I(\t0pre[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__A1 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3751__I (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3752__A1 (.I(\t0pre[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3753__A1 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3754__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3755__A1 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__A1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__C (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3757__A1 (.I(\t0pre[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3758__A1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__A1 (.I(\t0pre[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3760__A1 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3761__A1 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3762__I (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3763__C (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3766__A1 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__I (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3769__I (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3772__A1 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__A1 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3777__I (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__A1 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__A2 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3782__A1 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__A2 (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__A3 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__A1 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__I (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__A1 (.I(\t1pre[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__A1 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3793__A1 (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3794__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3795__A1 (.I(\t1pre[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3796__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__A1 (.I(\t1pre[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3799__A1 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3801__A1 (.I(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3802__A1 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3806__I (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3807__A1 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3808__A1 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3809__A1 (.I(\t1pre[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3810__A1 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3812__A1 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__C (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3815__A1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__A1 (.I(\t1pre[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3817__A1 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__A1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__I (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3823__I (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3825__A1 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3826__A1 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__A1 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__I (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3829__C (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3831__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3831__C (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3832__A1 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__C (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__A1 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__A2 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__A1 (.I(\t2pre[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__A3 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__I (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3840__A1 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3842__B (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3844__I (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__I (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__A1 (.I(\t2pre[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__A1 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3848__A1 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3849__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__A1 (.I(\t2pre[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3851__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__A1 (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3854__A1 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3855__B (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3856__A1 (.I(\t2pre[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3857__A1 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__I (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__I (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__A1 (.I(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3862__A1 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3863__A1 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__A1 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__A1 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__A1 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__C (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__A1 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__A1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__A1 (.I(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__A1 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__A1 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__C (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__A1 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__C (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__A1 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__I (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__C (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__C (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__A1 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__C (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__A2 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__A1 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__A2 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__A1 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3895__I (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3908__I (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3909__I (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3922__I (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3930__A2 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3932__I (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__A2 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3935__A2 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3937__I (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__A2 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__A1 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__A2 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__I (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__I (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__I (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__A1 (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__I (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__I (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3959__I (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3967__I (.I(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__I (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__I (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__I (.I(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__A2 (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__B1 (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__A1 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3994__A2 (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3994__B1 (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__A1 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__A2 (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__B1 (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__A1 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__I (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4003__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4003__A2 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4004__A1 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__A2 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4008__A2 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__A2 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4010__C (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__B (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__I (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4014__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4014__A2 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__A1 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4019__A1 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4019__A2 (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4019__C (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__I (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__A1 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__A1 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__C (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__A2 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__A4 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__A2 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A1 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__C (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4040__A2 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__A1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__A2 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__A1 (.I(\timer2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__I (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__A1 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__A1 (.I(\timer2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__A2 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4050__A1 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__A1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4053__I (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4054__A1 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4054__A2 (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4054__C (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__A1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__A1 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__I (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4060__A1 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__A2 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__A3 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__A2 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__A1 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__I (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__A1 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__A1 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__A2 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__A1 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__A1 (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__A2 (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__C (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4080__A1 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__A1 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__C (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4082__A1 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__A1 (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__A1 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__A1 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4089__A1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__B (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__A1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4094__B2 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4095__A1 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__A1 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__A1 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__A2 (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__C (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__A2 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4111__B2 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4112__A1 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4112__A2 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4112__B (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4114__A2 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4116__A1 (.I(\t0_top[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4117__A1 (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__I (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__A1 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__A1 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A1 (.I(\t0_top[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4124__A1 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4124__C (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__I (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4128__A1 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4129__I (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__A1 (.I(\t0_top[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__A1 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4136__A1 (.I(\temp[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A1 (.I(\temp[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__C (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__A1 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__C (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__A1 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__C (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4148__A1 (.I(\t0_top[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__A1 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__C (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A1 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4155__A1 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__A1 (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__A1 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4163__I (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A1 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__I (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4170__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4172__I (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4173__A1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4175__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4177__A1 (.I(\t1_top[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4178__A1 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4179__A1 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4182__A1 (.I(\t1_top[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__I (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__I (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4185__A1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4186__A1 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__A1 (.I(\temp[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4190__A1 (.I(\t1_top[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4191__A1 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4192__A1 (.I(\t1_top[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4193__I (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__A1 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__I (.I(\t1_top[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__A1 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__A1 (.I(\t1_top[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__A1 (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4201__A1 (.I(\t1_top[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__A1 (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__I (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__A1 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__I (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__A1 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4211__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4347__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4413__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__D (.I(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_wb_clk_i_I (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_wb_clk_i_I (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_wb_clk_i_I (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_wb_clk_i_I (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_wb_clk_i_I (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_wb_clk_i_I (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_wb_clk_i_I (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_wb_clk_i_I (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_wb_clk_i_I (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_wb_clk_i_I (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_wb_clk_i_I (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_wb_clk_i_I (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_wb_clk_i_I (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_wb_clk_i_I (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_wb_clk_i_I (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_wb_clk_i_I (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_wb_clk_i_I (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_wb_clk_i_I (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_wb_clk_i_I (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_wb_clk_i_I (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_wb_clk_i_I (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_wb_clk_i_I (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_wb_clk_i_I (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_64_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_70_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_72_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_73_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_78_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_81_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_82_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_83_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_84_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_85_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_86_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_87_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_88_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_89_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_90_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_91_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_92_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_93_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(data_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(data_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(data_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(data_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(data_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(data_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(data_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(rst));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(tmr0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(tmr1_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(bus_cyc));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(bus_we));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(data_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output20_I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output21_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output23_I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output24_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output28_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output29_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output31_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output32_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Left_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Left_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Left_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Left_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Left_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Left_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Left_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Left_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Left_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Left_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Left_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Left_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Left_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Left_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Left_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Left_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Left_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Left_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Left_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Left_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Left_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Left_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Left_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Left_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Left_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Left_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Left_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Left_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Left_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_310 ();
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2104_ (.A1(_0591_),
    .A2(_1638_),
    .B(_1645_),
    .C(_1644_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2105_ (.A1(_1320_),
    .A2(_1642_),
    .ZN(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2106_ (.A1(_0605_),
    .A2(_1638_),
    .B(_1646_),
    .C(_1644_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2107_ (.A1(_1322_),
    .A2(_1642_),
    .ZN(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2108_ (.A1(_0587_),
    .A2(_1619_),
    .B(_1647_),
    .C(_1644_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2109_ (.A1(_1614_),
    .A2(_1617_),
    .ZN(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2110_ (.I(_1630_),
    .Z(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2111_ (.A1(_0609_),
    .A2(_1619_),
    .B(_1648_),
    .C(_1649_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2112_ (.A1(_1869_),
    .A2(_1846_),
    .A3(_1278_),
    .ZN(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2113_ (.I(_1650_),
    .Z(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2114_ (.I(_1651_),
    .Z(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2115_ (.I(_1650_),
    .Z(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2116_ (.I(_1653_),
    .Z(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2117_ (.A1(_1056_),
    .A2(_1654_),
    .ZN(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2118_ (.A1(_0910_),
    .A2(_1652_),
    .B(_1655_),
    .C(_1649_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2119_ (.I(_1653_),
    .Z(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2120_ (.A1(_0962_),
    .A2(_1656_),
    .ZN(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2121_ (.A1(_0907_),
    .A2(_1652_),
    .B(_1657_),
    .C(_1649_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2122_ (.A1(\temp[2] ),
    .A2(_1656_),
    .ZN(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2123_ (.A1(_0903_),
    .A2(_1652_),
    .B(_1658_),
    .C(_1649_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2124_ (.A1(\temp[3] ),
    .A2(_1656_),
    .ZN(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2125_ (.I(_1356_),
    .Z(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2126_ (.A1(_0901_),
    .A2(_1652_),
    .B(_1659_),
    .C(_1660_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2127_ (.I(_1651_),
    .Z(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2128_ (.A1(_0989_),
    .A2(_1656_),
    .ZN(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2129_ (.A1(_0899_),
    .A2(_1661_),
    .B(_1662_),
    .C(_1660_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2130_ (.I(_1653_),
    .Z(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2131_ (.A1(\temp[5] ),
    .A2(_1663_),
    .ZN(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2132_ (.A1(_0897_),
    .A2(_1661_),
    .B(_1664_),
    .C(_1660_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2133_ (.A1(\temp[6] ),
    .A2(_1663_),
    .ZN(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2134_ (.A1(_0894_),
    .A2(_1661_),
    .B(_1665_),
    .C(_1660_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2135_ (.A1(_1008_),
    .A2(_1663_),
    .ZN(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2136_ (.I(_1356_),
    .Z(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2137_ (.A1(_0891_),
    .A2(_1661_),
    .B(_1666_),
    .C(_1667_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2138_ (.I(_1651_),
    .Z(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2139_ (.A1(_1308_),
    .A2(_1663_),
    .ZN(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2140_ (.A1(_0875_),
    .A2(_1668_),
    .B(_1669_),
    .C(_1667_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2141_ (.I(_1653_),
    .Z(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2142_ (.A1(net10),
    .A2(_1670_),
    .ZN(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2143_ (.A1(_0872_),
    .A2(_1668_),
    .B(_1671_),
    .C(_1667_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2144_ (.A1(net11),
    .A2(_1670_),
    .ZN(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2145_ (.A1(_0877_),
    .A2(_1668_),
    .B(_1672_),
    .C(_1667_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2146_ (.A1(_1028_),
    .A2(_1670_),
    .ZN(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2147_ (.I(_1356_),
    .Z(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2148_ (.A1(_0879_),
    .A2(_1668_),
    .B(_1673_),
    .C(_1674_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2149_ (.A1(_1875_),
    .A2(_0973_),
    .ZN(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2150_ (.A1(_1998_),
    .A2(_1675_),
    .ZN(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2151_ (.A1(_1039_),
    .A2(_1654_),
    .ZN(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2152_ (.A1(_0646_),
    .A2(_1676_),
    .A3(_1677_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2153_ (.A1(_2016_),
    .A2(_1675_),
    .ZN(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2154_ (.A1(_1041_),
    .A2(_1675_),
    .B(_1678_),
    .C(_1674_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2155_ (.A1(_1322_),
    .A2(_1670_),
    .ZN(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2156_ (.A1(_0887_),
    .A2(_1654_),
    .B(_1679_),
    .C(_1674_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2157_ (.A1(_1614_),
    .A2(_1651_),
    .ZN(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2158_ (.A1(_0863_),
    .A2(_1654_),
    .B(_1680_),
    .C(_1674_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2159_ (.A1(_0464_),
    .A2(_1485_),
    .ZN(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2160_ (.I(_1681_),
    .Z(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2161_ (.I(_1682_),
    .Z(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2162_ (.A1(_0828_),
    .A2(_1683_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2163_ (.A1(_0834_),
    .A2(_1683_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2164_ (.A1(_0830_),
    .A2(_1683_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2165_ (.A1(_0832_),
    .A2(_1683_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2166_ (.I(_1681_),
    .Z(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2167_ (.A1(_0821_),
    .A2(_1684_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2168_ (.A1(_0841_),
    .A2(_1684_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2169_ (.A1(_0826_),
    .A2(_1684_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2170_ (.A1(_0808_),
    .A2(_1684_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2171_ (.I(_1681_),
    .Z(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2172_ (.A1(_0801_),
    .A2(_1685_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2173_ (.A1(_0793_),
    .A2(_1685_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2174_ (.A1(_0786_),
    .A2(_1685_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2175_ (.A1(_0789_),
    .A2(_1685_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2176_ (.A1(_0468_),
    .A2(_0773_),
    .A3(_1502_),
    .Z(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2177_ (.I(_1686_),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2178_ (.A1(_0765_),
    .A2(_0764_),
    .A3(_1682_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2179_ (.A1(_0758_),
    .A2(_1682_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2180_ (.A1(_0762_),
    .A2(_1682_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2181_ (.A1(_0654_),
    .A2(_1782_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2182_ (.A1(_0654_),
    .A2(\pwm_ctr0[1] ),
    .ZN(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2183_ (.A1(_0740_),
    .A2(_1687_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2184_ (.I(_1788_),
    .Z(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2185_ (.I(_0668_),
    .Z(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2186_ (.A1(_0654_),
    .A2(\pwm_ctr0[1] ),
    .B(\pwm_ctr0[2] ),
    .ZN(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2187_ (.A1(_1688_),
    .A2(_1689_),
    .A3(_1690_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2188_ (.A1(_0657_),
    .A2(_1689_),
    .B(_1044_),
    .ZN(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2189_ (.A1(_0657_),
    .A2(_1689_),
    .B(_1691_),
    .ZN(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2190_ (.I(_1692_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2191_ (.A1(_0657_),
    .A2(_1689_),
    .B(\pwm_ctr0[4] ),
    .ZN(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2192_ (.A1(_1688_),
    .A2(_0669_),
    .A3(_1693_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2193_ (.A1(\pwm_ctr0[5] ),
    .A2(_0669_),
    .ZN(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2194_ (.A1(_1688_),
    .A2(_0670_),
    .A3(_1694_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2195_ (.A1(_0652_),
    .A2(_0670_),
    .ZN(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2196_ (.A1(_0652_),
    .A2(_0670_),
    .Z(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2197_ (.A1(_0946_),
    .A2(_1695_),
    .A3(_1696_),
    .ZN(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2198_ (.I(_1697_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2199_ (.A1(_0468_),
    .A2(_0671_),
    .ZN(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2200_ (.A1(_0659_),
    .A2(_1695_),
    .B(_1698_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2201_ (.A1(_0678_),
    .A2(_1782_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2202_ (.A1(_0678_),
    .A2(\pwm_ctr1[1] ),
    .ZN(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2203_ (.A1(_0740_),
    .A2(_1699_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2204_ (.I(_0692_),
    .Z(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2205_ (.A1(_0678_),
    .A2(\pwm_ctr1[1] ),
    .B(\pwm_ctr1[2] ),
    .ZN(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2206_ (.A1(_1688_),
    .A2(_1700_),
    .A3(_1701_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2207_ (.A1(_0681_),
    .A2(_1700_),
    .B(_1044_),
    .ZN(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2208_ (.A1(_0681_),
    .A2(_1700_),
    .B(_1702_),
    .ZN(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2209_ (.I(_1703_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2210_ (.A1(_0681_),
    .A2(_1700_),
    .B(\pwm_ctr1[4] ),
    .ZN(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2211_ (.A1(_0988_),
    .A2(_0693_),
    .A3(_1704_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2212_ (.A1(\pwm_ctr1[5] ),
    .A2(_0693_),
    .ZN(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2213_ (.A1(_0988_),
    .A2(_0694_),
    .A3(_1705_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2214_ (.A1(_0676_),
    .A2(_0694_),
    .ZN(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2215_ (.A1(_0676_),
    .A2(_0694_),
    .Z(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2216_ (.A1(_0946_),
    .A2(_1706_),
    .A3(_1707_),
    .ZN(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2217_ (.I(_1708_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2218_ (.A1(_0468_),
    .A2(_0695_),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2219_ (.A1(_0683_),
    .A2(_1706_),
    .B(_1709_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2220_ (.A1(_1989_),
    .A2(_0973_),
    .ZN(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2221_ (.A1(\pw0[0] ),
    .A2(_1710_),
    .ZN(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2222_ (.A1(_1879_),
    .A2(_0719_),
    .Z(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2223_ (.I(_1712_),
    .Z(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2224_ (.A1(_0724_),
    .A2(_1713_),
    .ZN(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2225_ (.A1(_1711_),
    .A2(_1714_),
    .B(_1371_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2226_ (.I(_1712_),
    .Z(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2227_ (.I(_1712_),
    .Z(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2228_ (.I(_1345_),
    .Z(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2229_ (.A1(\pw0[1] ),
    .A2(_1716_),
    .B(_1717_),
    .ZN(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2230_ (.A1(_1604_),
    .A2(_1715_),
    .B(_1718_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2231_ (.I(_0731_),
    .Z(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2232_ (.A1(\pw0[2] ),
    .A2(_1716_),
    .B(_1717_),
    .ZN(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2233_ (.A1(_1719_),
    .A2(_1715_),
    .B(_1720_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2234_ (.A1(\pw0[3] ),
    .A2(_1710_),
    .ZN(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2235_ (.A1(_1354_),
    .A2(_1713_),
    .ZN(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2236_ (.I(_1245_),
    .Z(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2237_ (.A1(_1721_),
    .A2(_1722_),
    .B(_1723_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2238_ (.A1(_0469_),
    .A2(_1710_),
    .ZN(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2239_ (.A1(_0651_),
    .A2(_1710_),
    .B(_1724_),
    .C(_1530_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2240_ (.A1(\pw0[5] ),
    .A2(_1716_),
    .B(_1717_),
    .ZN(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2241_ (.A1(_1610_),
    .A2(_1715_),
    .B(_1725_),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2242_ (.A1(\pw0[6] ),
    .A2(_1716_),
    .B(_1717_),
    .ZN(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2243_ (.A1(_0736_),
    .A2(_1715_),
    .B(_1726_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2244_ (.A1(_1614_),
    .A2(_1713_),
    .ZN(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2245_ (.A1(_0661_),
    .A2(_1713_),
    .B(_1727_),
    .C(_1357_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2246_ (.A1(_1905_),
    .A2(_0973_),
    .ZN(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2247_ (.A1(\pw1[0] ),
    .A2(_1728_),
    .ZN(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2248_ (.A1(_1841_),
    .A2(_1878_),
    .A3(_0460_),
    .ZN(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2249_ (.I(_1730_),
    .Z(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2250_ (.A1(_1546_),
    .A2(_1731_),
    .ZN(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2251_ (.A1(_1729_),
    .A2(_1732_),
    .B(_1723_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2252_ (.I(_1730_),
    .Z(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2253_ (.I(_1730_),
    .Z(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2254_ (.I(_1317_),
    .Z(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2255_ (.A1(\pw1[1] ),
    .A2(_1734_),
    .B(_1735_),
    .ZN(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2256_ (.A1(_1604_),
    .A2(_1733_),
    .B(_1736_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2257_ (.A1(\pw1[2] ),
    .A2(_1734_),
    .B(_1735_),
    .ZN(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2258_ (.A1(_1719_),
    .A2(_1733_),
    .B(_1737_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2259_ (.A1(\pw1[3] ),
    .A2(_1728_),
    .ZN(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2260_ (.A1(_1354_),
    .A2(_1731_),
    .ZN(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2261_ (.A1(_1738_),
    .A2(_1739_),
    .B(_1723_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2262_ (.A1(_1038_),
    .A2(_1728_),
    .ZN(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2263_ (.I(_0987_),
    .Z(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2264_ (.A1(_0675_),
    .A2(_1728_),
    .B(_1740_),
    .C(_1741_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2265_ (.A1(\pw1[5] ),
    .A2(_1734_),
    .B(_1735_),
    .ZN(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2266_ (.A1(_1610_),
    .A2(_1733_),
    .B(_1742_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2267_ (.A1(\pw1[6] ),
    .A2(_1734_),
    .B(_1735_),
    .ZN(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2268_ (.A1(_0736_),
    .A2(_1733_),
    .B(_1743_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2269_ (.A1(_1052_),
    .A2(_1731_),
    .ZN(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2270_ (.A1(_0685_),
    .A2(_1731_),
    .B(_1744_),
    .C(_1357_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2271_ (.A1(_1881_),
    .A2(_1273_),
    .ZN(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2272_ (.I(_1745_),
    .Z(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2273_ (.A1(_0723_),
    .A2(_1746_),
    .ZN(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2274_ (.A1(_0697_),
    .A2(_1746_),
    .B(_1747_),
    .C(_1741_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2275_ (.A1(_1878_),
    .A2(_1853_),
    .A3(_1278_),
    .ZN(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2276_ (.I(_1748_),
    .Z(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2277_ (.I(_1748_),
    .Z(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2278_ (.I(_1317_),
    .Z(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2279_ (.A1(\pw2[1] ),
    .A2(_1750_),
    .B(_1751_),
    .ZN(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2280_ (.A1(_1604_),
    .A2(_1749_),
    .B(_1752_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2281_ (.A1(\pw2[2] ),
    .A2(_1750_),
    .B(_1751_),
    .ZN(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2282_ (.A1(_1719_),
    .A2(_1749_),
    .B(_1753_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2283_ (.A1(_1142_),
    .A2(_1745_),
    .ZN(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2284_ (.A1(_0706_),
    .A2(_1746_),
    .B(_1754_),
    .C(_1741_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2285_ (.A1(_1038_),
    .A2(_1745_),
    .ZN(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2286_ (.A1(_0702_),
    .A2(_1746_),
    .B(_1755_),
    .C(_1741_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2287_ (.A1(\pw2[5] ),
    .A2(_1748_),
    .B(_1751_),
    .ZN(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2288_ (.A1(_1610_),
    .A2(_1749_),
    .B(_1756_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2289_ (.A1(\pw2[6] ),
    .A2(_1748_),
    .B(_1751_),
    .ZN(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2290_ (.A1(_0736_),
    .A2(_1749_),
    .B(_1757_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2291_ (.A1(_1052_),
    .A2(_1750_),
    .ZN(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2292_ (.A1(_0707_),
    .A2(_1750_),
    .B(_1758_),
    .C(_1357_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2293_ (.A1(_1808_),
    .A2(_1814_),
    .B(_1825_),
    .ZN(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2294_ (.A1(_1854_),
    .A2(_1759_),
    .B(_1810_),
    .ZN(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2295_ (.A1(_1893_),
    .A2(_1760_),
    .B(_0718_),
    .ZN(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2296_ (.I(_1761_),
    .Z(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2297_ (.A1(\temp[0] ),
    .A2(_1762_),
    .ZN(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2298_ (.A1(_1894_),
    .A2(_1760_),
    .ZN(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2299_ (.A1(_0460_),
    .A2(_1764_),
    .ZN(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2300_ (.A1(_1546_),
    .A2(_1765_),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2301_ (.A1(_1763_),
    .A2(_1766_),
    .B(_1723_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2302_ (.I(_1761_),
    .Z(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2303_ (.A1(net10),
    .A2(_1762_),
    .ZN(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2304_ (.I(_0987_),
    .Z(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2305_ (.A1(_1283_),
    .A2(_1767_),
    .B(_1768_),
    .C(_1769_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2306_ (.A1(\temp[2] ),
    .A2(_1765_),
    .B(_1318_),
    .ZN(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2307_ (.A1(_1719_),
    .A2(_1765_),
    .B(_1770_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2308_ (.I(_1761_),
    .Z(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2309_ (.A1(_0457_),
    .A2(_1771_),
    .ZN(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2310_ (.A1(_0980_),
    .A2(_1767_),
    .B(_1772_),
    .C(_1769_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2311_ (.A1(\temp[4] ),
    .A2(_1762_),
    .ZN(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2312_ (.A1(_1315_),
    .A2(_1765_),
    .ZN(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2313_ (.A1(_1773_),
    .A2(_1774_),
    .B(_1785_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2314_ (.A1(_0717_),
    .A2(_1771_),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2315_ (.A1(_0997_),
    .A2(_1767_),
    .B(_1775_),
    .C(_1769_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2316_ (.A1(net15),
    .A2(_1771_),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2317_ (.A1(_1001_),
    .A2(_1767_),
    .B(_1776_),
    .C(_1769_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2318_ (.A1(_0738_),
    .A2(_1771_),
    .ZN(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2319_ (.A1(_1305_),
    .A2(_1762_),
    .B(_1777_),
    .C(_1789_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2320_ (.I(\pwm_ctr2[0] ),
    .Z(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2321_ (.I(net17),
    .Z(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2322_ (.I(_1779_),
    .Z(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2323_ (.I(_1780_),
    .Z(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2324_ (.I(_1781_),
    .Z(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2325_ (.A1(_1778_),
    .A2(_1782_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2326_ (.I(net17),
    .Z(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2327_ (.I(_1783_),
    .Z(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2328_ (.I(_1784_),
    .Z(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2329_ (.I(\pwm_ctr2[1] ),
    .ZN(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2330_ (.A1(_1778_),
    .A2(_1786_),
    .Z(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2331_ (.A1(_1785_),
    .A2(_1787_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2332_ (.I(_1779_),
    .Z(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2333_ (.I(_1788_),
    .Z(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2334_ (.A1(_1778_),
    .A2(\pwm_ctr2[1] ),
    .B(\pwm_ctr2[2] ),
    .ZN(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2335_ (.A1(\pwm_ctr2[0] ),
    .A2(\pwm_ctr2[1] ),
    .A3(\pwm_ctr2[2] ),
    .Z(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2336_ (.A1(_1789_),
    .A2(_1790_),
    .A3(_1791_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2337_ (.A1(\pwm_ctr2[3] ),
    .A2(_1791_),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2338_ (.A1(\pwm_ctr2[3] ),
    .A2(_1791_),
    .Z(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2339_ (.A1(_1789_),
    .A2(_1792_),
    .A3(_1793_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2340_ (.A1(\pwm_ctr2[4] ),
    .A2(_1793_),
    .ZN(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2341_ (.A1(\pwm_ctr2[4] ),
    .A2(_1793_),
    .Z(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2342_ (.A1(_1789_),
    .A2(_1794_),
    .A3(_1795_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2343_ (.I(_1788_),
    .Z(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2344_ (.A1(\pwm_ctr2[5] ),
    .A2(_1795_),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2345_ (.A1(\pwm_ctr2[5] ),
    .A2(_1795_),
    .Z(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2346_ (.A1(_1796_),
    .A2(_1797_),
    .A3(_1798_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2347_ (.A1(\pwm_ctr2[6] ),
    .A2(_1798_),
    .ZN(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2348_ (.A1(\pwm_ctr2[6] ),
    .A2(_1798_),
    .Z(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2349_ (.A1(_1796_),
    .A2(_1799_),
    .A3(_1800_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2350_ (.I(\pwm_ctr2[7] ),
    .Z(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2351_ (.I(net17),
    .ZN(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2352_ (.I(_1802_),
    .Z(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2353_ (.I(_1803_),
    .Z(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2354_ (.I(_1804_),
    .Z(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2355_ (.A1(_1801_),
    .A2(_1800_),
    .B(_1805_),
    .ZN(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2356_ (.A1(_1801_),
    .A2(_1800_),
    .B(_1806_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2357_ (.I(net2),
    .Z(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2358_ (.I(_1807_),
    .Z(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2359_ (.I(net1),
    .Z(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2360_ (.I(_1809_),
    .Z(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2361_ (.I(net5),
    .ZN(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2362_ (.A1(net6),
    .A2(_1811_),
    .ZN(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2363_ (.I(net3),
    .Z(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2364_ (.I(net4),
    .Z(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2365_ (.A1(_1813_),
    .A2(_1814_),
    .ZN(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2366_ (.A1(_1812_),
    .A2(_1815_),
    .ZN(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2367_ (.A1(_1808_),
    .A2(_1810_),
    .A3(_1816_),
    .ZN(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2368_ (.I(_1817_),
    .Z(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2369_ (.I(net3),
    .ZN(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2370_ (.I(net4),
    .ZN(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2371_ (.A1(_1819_),
    .A2(_1820_),
    .ZN(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2372_ (.I(_1821_),
    .Z(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2373_ (.I(net1),
    .ZN(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2374_ (.A1(net6),
    .A2(net5),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2375_ (.I(_1824_),
    .Z(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2376_ (.A1(_1807_),
    .A2(_1823_),
    .A3(_1825_),
    .ZN(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2377_ (.A1(_1822_),
    .A2(_1826_),
    .ZN(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2378_ (.I(_1827_),
    .Z(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2379_ (.A1(\t1_capture[0] ),
    .A2(_1818_),
    .B1(_1828_),
    .B2(\t0pre[0] ),
    .ZN(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2380_ (.A1(_1807_),
    .A2(_1809_),
    .A3(_1824_),
    .ZN(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2381_ (.I(_1830_),
    .Z(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2382_ (.A1(_1831_),
    .A2(_1821_),
    .ZN(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2383_ (.I(_1832_),
    .Z(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2384_ (.I(net2),
    .ZN(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2385_ (.A1(_1834_),
    .A2(_1823_),
    .A3(_1825_),
    .ZN(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2386_ (.A1(_1821_),
    .A2(_1835_),
    .ZN(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2387_ (.I(_1836_),
    .Z(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2388_ (.I(_1837_),
    .Z(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2389_ (.A1(\t0pre[8] ),
    .A2(_1833_),
    .B1(_1838_),
    .B2(\settings[0] ),
    .ZN(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2390_ (.A1(_1834_),
    .A2(_1809_),
    .ZN(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2391_ (.I(_1840_),
    .Z(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2392_ (.A1(_1841_),
    .A2(_1816_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2393_ (.I(_1842_),
    .Z(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2394_ (.I(_1835_),
    .Z(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2395_ (.A1(_1813_),
    .A2(_1814_),
    .ZN(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2396_ (.I(_1845_),
    .Z(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2397_ (.A1(_1844_),
    .A2(_1846_),
    .ZN(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2398_ (.I(_1847_),
    .Z(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2399_ (.A1(\t1_capture[8] ),
    .A2(_1843_),
    .B1(_1848_),
    .B2(\t2_top[0] ),
    .ZN(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2400_ (.A1(_1813_),
    .A2(_1820_),
    .ZN(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2401_ (.A1(_1850_),
    .A2(_1831_),
    .ZN(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2402_ (.I(_1851_),
    .Z(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2403_ (.A1(_1808_),
    .A2(_1823_),
    .ZN(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2404_ (.I(_1816_),
    .Z(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2405_ (.A1(_1853_),
    .A2(_1854_),
    .ZN(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2406_ (.I(_1855_),
    .Z(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2407_ (.A1(\t2pre[8] ),
    .A2(_1852_),
    .B1(_1856_),
    .B2(\t2_capture[0] ),
    .ZN(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2408_ (.A1(_1829_),
    .A2(_1839_),
    .A3(_1849_),
    .A4(_1857_),
    .ZN(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2409_ (.A1(_1834_),
    .A2(_1809_),
    .A3(_1825_),
    .ZN(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2410_ (.A1(_1819_),
    .A2(_1814_),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2411_ (.A1(_1859_),
    .A2(_1860_),
    .ZN(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2412_ (.I(_1861_),
    .Z(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2413_ (.A1(\t0_top[8] ),
    .A2(_1862_),
    .ZN(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2414_ (.A1(net6),
    .A2(net5),
    .A3(_1840_),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2415_ (.I(net7),
    .ZN(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2416_ (.A1(_1864_),
    .A2(_1815_),
    .B(net17),
    .C(_1865_),
    .ZN(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2417_ (.I(_1866_),
    .Z(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2418_ (.I(_1850_),
    .Z(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2419_ (.I(_1859_),
    .Z(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2420_ (.A1(_1868_),
    .A2(_1869_),
    .ZN(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2421_ (.I(_1870_),
    .Z(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2422_ (.A1(_1826_),
    .A2(_1846_),
    .ZN(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2423_ (.I(_1872_),
    .Z(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2424_ (.A1(_1859_),
    .A2(_1845_),
    .ZN(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2425_ (.I(_1874_),
    .Z(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _2426_ (.A1(\t1pre[8] ),
    .A2(_1871_),
    .B1(_1873_),
    .B2(\t0_capture[0] ),
    .C1(_1875_),
    .C2(\t2_top[8] ),
    .ZN(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2427_ (.A1(_1813_),
    .A2(_1820_),
    .A3(_1812_),
    .ZN(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2428_ (.I(_1877_),
    .Z(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2429_ (.A1(_1808_),
    .A2(_1810_),
    .A3(_1878_),
    .ZN(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2430_ (.A1(_1877_),
    .A2(_1853_),
    .ZN(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2431_ (.I(_1880_),
    .Z(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2432_ (.A1(\pw0[0] ),
    .A2(_1879_),
    .B1(_1881_),
    .B2(\pw2[0] ),
    .ZN(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2433_ (.A1(_1863_),
    .A2(_1867_),
    .A3(_1876_),
    .A4(_1882_),
    .ZN(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2434_ (.I(_1860_),
    .Z(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2435_ (.A1(_1884_),
    .A2(_1844_),
    .ZN(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2436_ (.I(_1885_),
    .Z(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2437_ (.A1(_1884_),
    .A2(_1826_),
    .ZN(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2438_ (.I(_1887_),
    .Z(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2439_ (.A1(\t0_top[0] ),
    .A2(_1886_),
    .B1(_1888_),
    .B2(\t1_top[0] ),
    .ZN(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2440_ (.A1(_1807_),
    .A2(_1810_),
    .ZN(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2441_ (.A1(_1890_),
    .A2(_1816_),
    .ZN(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2442_ (.I(_1891_),
    .Z(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2443_ (.A1(_1868_),
    .A2(_1844_),
    .ZN(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2444_ (.I(_1893_),
    .Z(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2445_ (.I(\t1pre[0] ),
    .Z(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2446_ (.A1(\t2_capture[8] ),
    .A2(_1892_),
    .B1(_1894_),
    .B2(_1895_),
    .ZN(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2447_ (.A1(_1831_),
    .A2(_1845_),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2448_ (.I(_1897_),
    .Z(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2449_ (.A1(_1850_),
    .A2(_1826_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2450_ (.I(_1899_),
    .Z(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2451_ (.A1(\t0_capture[8] ),
    .A2(_1898_),
    .B1(_1900_),
    .B2(\t2pre[0] ),
    .ZN(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2452_ (.A1(_1831_),
    .A2(_1860_),
    .ZN(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2453_ (.I(_1902_),
    .Z(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2454_ (.A1(_1841_),
    .A2(_1878_),
    .ZN(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2455_ (.I(_1904_),
    .Z(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2456_ (.A1(\t1_top[8] ),
    .A2(_1903_),
    .B1(_1905_),
    .B2(\pw1[0] ),
    .ZN(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2457_ (.A1(_1889_),
    .A2(_1896_),
    .A3(_1901_),
    .A4(_1906_),
    .ZN(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2458_ (.A1(_1783_),
    .A2(_1865_),
    .ZN(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2459_ (.I(_1908_),
    .Z(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2460_ (.A1(_1858_),
    .A2(_1883_),
    .A3(_1907_),
    .B1(_1909_),
    .B2(net20),
    .ZN(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2461_ (.I(_1910_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2462_ (.I(_1908_),
    .Z(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2463_ (.I(_1902_),
    .Z(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2464_ (.I(_1899_),
    .Z(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2465_ (.A1(\t1_top[9] ),
    .A2(_1912_),
    .B1(_1913_),
    .B2(\t2pre[1] ),
    .ZN(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2466_ (.I(_1885_),
    .Z(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2467_ (.I(_1855_),
    .Z(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2468_ (.A1(\t0_top[1] ),
    .A2(_1915_),
    .B1(_1916_),
    .B2(\t2_capture[1] ),
    .ZN(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2469_ (.I(_1817_),
    .Z(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2470_ (.I(_1827_),
    .Z(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2471_ (.A1(\t1_capture[1] ),
    .A2(_1918_),
    .B1(_1919_),
    .B2(\t0pre[1] ),
    .ZN(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2472_ (.I(_1879_),
    .Z(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2473_ (.I(_1851_),
    .Z(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2474_ (.I(\t2pre[9] ),
    .Z(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2475_ (.A1(\pw0[1] ),
    .A2(_1921_),
    .B1(_1922_),
    .B2(_1923_),
    .ZN(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2476_ (.A1(_1914_),
    .A2(_1917_),
    .A3(_1920_),
    .A4(_1924_),
    .ZN(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2477_ (.I(_1880_),
    .Z(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2478_ (.I(_1842_),
    .Z(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2479_ (.A1(\pw2[1] ),
    .A2(_1926_),
    .B1(_1927_),
    .B2(\t1_capture[9] ),
    .ZN(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2480_ (.I(\t1pre[9] ),
    .Z(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2481_ (.I(_1870_),
    .Z(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2482_ (.I(_1893_),
    .Z(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2483_ (.A1(_1929_),
    .A2(_1930_),
    .B1(_1931_),
    .B2(\t1pre[1] ),
    .ZN(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2484_ (.I(_1872_),
    .Z(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _2485_ (.A1(\t2_top[1] ),
    .A2(_1848_),
    .B1(_1933_),
    .B2(\t0_capture[1] ),
    .C1(_1838_),
    .C2(\settings[1] ),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2486_ (.A1(\t0_capture[9] ),
    .A2(_1898_),
    .ZN(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2487_ (.A1(\t0_top[9] ),
    .A2(_1862_),
    .B1(_1875_),
    .B2(\t2_top[9] ),
    .ZN(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2488_ (.A1(\t0pre[9] ),
    .A2(_1833_),
    .B1(_1892_),
    .B2(\t2_capture[9] ),
    .ZN(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2489_ (.A1(_1867_),
    .A2(_1935_),
    .A3(_1936_),
    .A4(_1937_),
    .ZN(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2490_ (.A1(\pw1[1] ),
    .A2(_1905_),
    .B1(_1888_),
    .B2(\t1_top[1] ),
    .C(_1938_),
    .ZN(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2491_ (.A1(_1928_),
    .A2(_1932_),
    .A3(_1934_),
    .A4(_1939_),
    .ZN(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2492_ (.A1(net21),
    .A2(_1911_),
    .B1(_1925_),
    .B2(_1940_),
    .ZN(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2493_ (.I(_1941_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2494_ (.I(\t2pre[2] ),
    .Z(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2495_ (.A1(\t1_top[10] ),
    .A2(_1912_),
    .B1(_1913_),
    .B2(_1942_),
    .ZN(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2496_ (.A1(\t0_top[2] ),
    .A2(_1915_),
    .B1(_1916_),
    .B2(\t2_capture[2] ),
    .ZN(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2497_ (.I(\t0pre[2] ),
    .Z(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2498_ (.A1(\t1_capture[2] ),
    .A2(_1918_),
    .B1(_1919_),
    .B2(_1945_),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2499_ (.I(\t2pre[10] ),
    .Z(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2500_ (.A1(\pw0[2] ),
    .A2(_1921_),
    .B1(_1922_),
    .B2(_1947_),
    .ZN(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2501_ (.A1(_1943_),
    .A2(_1944_),
    .A3(_1946_),
    .A4(_1948_),
    .ZN(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2502_ (.A1(\pw2[2] ),
    .A2(_1926_),
    .B1(_1927_),
    .B2(\t1_capture[10] ),
    .ZN(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2503_ (.I(\t1pre[2] ),
    .Z(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2504_ (.A1(\t1pre[10] ),
    .A2(_1930_),
    .B1(_1931_),
    .B2(_1951_),
    .ZN(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _2505_ (.A1(\t2_top[2] ),
    .A2(_1848_),
    .B1(_1933_),
    .B2(\t0_capture[2] ),
    .C1(_1838_),
    .C2(\settings[2] ),
    .ZN(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2506_ (.I(_1897_),
    .Z(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2507_ (.A1(\t0_capture[10] ),
    .A2(_1954_),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2508_ (.I(_1861_),
    .Z(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2509_ (.I(_1874_),
    .Z(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2510_ (.A1(\t0_top[10] ),
    .A2(_1956_),
    .B1(_1957_),
    .B2(\t2_top[10] ),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2511_ (.I(_1832_),
    .Z(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2512_ (.I(_1891_),
    .Z(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2513_ (.A1(\t0pre[10] ),
    .A2(_1959_),
    .B1(_1960_),
    .B2(\t2_capture[10] ),
    .ZN(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2514_ (.A1(_1867_),
    .A2(_1955_),
    .A3(_1958_),
    .A4(_1961_),
    .ZN(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2515_ (.A1(\pw1[2] ),
    .A2(_1905_),
    .B1(_1888_),
    .B2(\t1_top[2] ),
    .C(_1962_),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2516_ (.A1(_1950_),
    .A2(_1952_),
    .A3(_1953_),
    .A4(_1963_),
    .ZN(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2517_ (.A1(net22),
    .A2(_1911_),
    .B1(_1949_),
    .B2(_1964_),
    .ZN(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2518_ (.I(_1965_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2519_ (.A1(\t1_top[11] ),
    .A2(_1912_),
    .B1(_1913_),
    .B2(\t2pre[3] ),
    .ZN(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2520_ (.A1(\t0_top[3] ),
    .A2(_1915_),
    .B1(_1916_),
    .B2(\t2_capture[3] ),
    .ZN(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2521_ (.A1(\t1_capture[3] ),
    .A2(_1918_),
    .B1(_1919_),
    .B2(\t0pre[3] ),
    .ZN(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2522_ (.A1(\pw0[3] ),
    .A2(_1921_),
    .B1(_1922_),
    .B2(\t2pre[11] ),
    .ZN(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2523_ (.A1(_1966_),
    .A2(_1967_),
    .A3(_1968_),
    .A4(_1969_),
    .ZN(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2524_ (.A1(\pw2[3] ),
    .A2(_1926_),
    .B1(_1927_),
    .B2(\t1_capture[11] ),
    .ZN(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2525_ (.I(\t1pre[11] ),
    .Z(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2526_ (.A1(_1972_),
    .A2(_1930_),
    .B1(_1931_),
    .B2(\t1pre[3] ),
    .ZN(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _2527_ (.A1(\t2_top[3] ),
    .A2(_1848_),
    .B1(_1933_),
    .B2(\t0_capture[3] ),
    .C1(_1838_),
    .C2(net28),
    .ZN(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2528_ (.I(_1904_),
    .Z(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2529_ (.I(_1866_),
    .Z(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2530_ (.A1(\t0_capture[11] ),
    .A2(_1954_),
    .ZN(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2531_ (.A1(\t0_top[11] ),
    .A2(_1956_),
    .B1(_1957_),
    .B2(\t2_top[11] ),
    .ZN(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2532_ (.A1(\t0pre[11] ),
    .A2(_1959_),
    .B1(_1960_),
    .B2(\t2_capture[11] ),
    .ZN(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2533_ (.A1(_1976_),
    .A2(_1977_),
    .A3(_1978_),
    .A4(_1979_),
    .ZN(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2534_ (.A1(\pw1[3] ),
    .A2(_1975_),
    .B1(_1888_),
    .B2(\t1_top[3] ),
    .C(_1980_),
    .ZN(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2535_ (.A1(_1971_),
    .A2(_1973_),
    .A3(_1974_),
    .A4(_1981_),
    .ZN(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2536_ (.A1(net23),
    .A2(_1911_),
    .B1(_1970_),
    .B2(_1982_),
    .ZN(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2537_ (.I(_1983_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2538_ (.I(\t2pre[4] ),
    .Z(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2539_ (.A1(\t1_top[12] ),
    .A2(_1912_),
    .B1(_1913_),
    .B2(_1984_),
    .ZN(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2540_ (.A1(\t0_top[4] ),
    .A2(_1915_),
    .B1(_1856_),
    .B2(\t2_capture[4] ),
    .ZN(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2541_ (.I(\t0pre[4] ),
    .Z(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2542_ (.A1(\t1_capture[4] ),
    .A2(_1918_),
    .B1(_1828_),
    .B2(_1987_),
    .ZN(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2543_ (.I(_1879_),
    .Z(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2544_ (.A1(\pw0[4] ),
    .A2(_1989_),
    .B1(_1922_),
    .B2(\t2pre[12] ),
    .ZN(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2545_ (.A1(_1985_),
    .A2(_1986_),
    .A3(_1988_),
    .A4(_1990_),
    .ZN(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2546_ (.A1(\pw2[4] ),
    .A2(_1926_),
    .B1(_1927_),
    .B2(\t1_capture[12] ),
    .ZN(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2547_ (.A1(\t1pre[12] ),
    .A2(_1930_),
    .B1(_1931_),
    .B2(\t1pre[4] ),
    .ZN(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2548_ (.I(_1847_),
    .Z(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _2549_ (.A1(\t2_top[4] ),
    .A2(_1994_),
    .B1(_1933_),
    .B2(\t0_capture[4] ),
    .C1(_1837_),
    .C2(net29),
    .ZN(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2550_ (.I(_1887_),
    .Z(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2551_ (.A1(\t0_capture[12] ),
    .A2(_1954_),
    .ZN(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2552_ (.I(\t2_top[12] ),
    .Z(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2553_ (.A1(\t0_top[12] ),
    .A2(_1956_),
    .B1(_1957_),
    .B2(_1998_),
    .ZN(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2554_ (.A1(\t0pre[12] ),
    .A2(_1959_),
    .B1(_1960_),
    .B2(\t2_capture[12] ),
    .ZN(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2555_ (.A1(_1976_),
    .A2(_1997_),
    .A3(_1999_),
    .A4(_2000_),
    .ZN(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2556_ (.A1(\pw1[4] ),
    .A2(_1975_),
    .B1(_1996_),
    .B2(\t1_top[4] ),
    .C(_2001_),
    .ZN(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2557_ (.A1(_1992_),
    .A2(_1993_),
    .A3(_1995_),
    .A4(_2002_),
    .ZN(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2558_ (.A1(net24),
    .A2(_1909_),
    .B1(_1991_),
    .B2(_2003_),
    .ZN(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2559_ (.I(_2004_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2560_ (.A1(\t1_top[13] ),
    .A2(_1903_),
    .B1(_1900_),
    .B2(\t2pre[5] ),
    .ZN(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2561_ (.A1(\t0_top[5] ),
    .A2(_1886_),
    .B1(_1856_),
    .B2(\t2_capture[5] ),
    .ZN(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2562_ (.I(\t0pre[5] ),
    .Z(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2563_ (.A1(\t1_capture[5] ),
    .A2(_1818_),
    .B1(_1828_),
    .B2(_2007_),
    .ZN(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2564_ (.A1(\pw0[5] ),
    .A2(_1989_),
    .B1(_1852_),
    .B2(\t2pre[13] ),
    .ZN(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2565_ (.A1(_2005_),
    .A2(_2006_),
    .A3(_2008_),
    .A4(_2009_),
    .ZN(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2566_ (.A1(\pw2[5] ),
    .A2(_1881_),
    .B1(_1843_),
    .B2(\t1_capture[13] ),
    .ZN(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2567_ (.I(\t1pre[5] ),
    .Z(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2568_ (.A1(\t1pre[13] ),
    .A2(_1871_),
    .B1(_1894_),
    .B2(_2012_),
    .ZN(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _2569_ (.A1(\t2_top[5] ),
    .A2(_1994_),
    .B1(_1873_),
    .B2(\t0_capture[5] ),
    .C1(_1837_),
    .C2(tmr0_ext),
    .ZN(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2570_ (.A1(\t0_capture[13] ),
    .A2(_1954_),
    .ZN(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2571_ (.I(\t2_top[13] ),
    .Z(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2572_ (.A1(\t0_top[13] ),
    .A2(_1956_),
    .B1(_1957_),
    .B2(_2016_),
    .ZN(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2573_ (.A1(\t0pre[13] ),
    .A2(_1959_),
    .B1(_1960_),
    .B2(\t2_capture[13] ),
    .ZN(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2574_ (.A1(_1976_),
    .A2(_2015_),
    .A3(_2017_),
    .A4(_2018_),
    .ZN(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2575_ (.A1(\pw1[5] ),
    .A2(_1975_),
    .B1(_1996_),
    .B2(\t1_top[5] ),
    .C(_2019_),
    .ZN(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2576_ (.A1(_2011_),
    .A2(_2013_),
    .A3(_2014_),
    .A4(_2020_),
    .ZN(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2577_ (.A1(net25),
    .A2(_1909_),
    .B1(_2010_),
    .B2(_2021_),
    .ZN(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2578_ (.I(_2022_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2579_ (.I(\t2pre[6] ),
    .Z(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2580_ (.A1(\t1_top[14] ),
    .A2(_1903_),
    .B1(_1900_),
    .B2(_2023_),
    .ZN(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2581_ (.A1(\t0_top[6] ),
    .A2(_1886_),
    .B1(_1856_),
    .B2(\t2_capture[6] ),
    .ZN(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2582_ (.A1(\t1_capture[6] ),
    .A2(_1818_),
    .B1(_1828_),
    .B2(\t0pre[6] ),
    .ZN(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2583_ (.A1(\pw0[6] ),
    .A2(_1989_),
    .B1(_1852_),
    .B2(\t2pre[14] ),
    .ZN(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2584_ (.A1(_2024_),
    .A2(_2025_),
    .A3(_2026_),
    .A4(_2027_),
    .ZN(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2585_ (.A1(\pw2[6] ),
    .A2(_1881_),
    .B1(_1843_),
    .B2(\t1_capture[14] ),
    .ZN(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2586_ (.I(\t1pre[6] ),
    .Z(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2587_ (.A1(\t1pre[14] ),
    .A2(_1871_),
    .B1(_1894_),
    .B2(_2030_),
    .ZN(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _2588_ (.A1(\t2_top[6] ),
    .A2(_1994_),
    .B1(_1873_),
    .B2(\t0_capture[6] ),
    .C1(_1837_),
    .C2(tmr1_ext),
    .ZN(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2589_ (.A1(\t0_capture[14] ),
    .A2(_1897_),
    .ZN(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2590_ (.A1(\t0_top[14] ),
    .A2(_1861_),
    .B1(_1874_),
    .B2(\t2_top[14] ),
    .ZN(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2591_ (.A1(\t0pre[14] ),
    .A2(_1832_),
    .B1(_1891_),
    .B2(\t2_capture[14] ),
    .ZN(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2592_ (.A1(_1976_),
    .A2(_2033_),
    .A3(_2034_),
    .A4(_2035_),
    .ZN(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2593_ (.A1(\pw1[6] ),
    .A2(_1975_),
    .B1(_1996_),
    .B2(\t1_top[6] ),
    .C(_2036_),
    .ZN(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2594_ (.A1(_2029_),
    .A2(_2031_),
    .A3(_2032_),
    .A4(_2037_),
    .ZN(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2595_ (.A1(net26),
    .A2(_1909_),
    .B1(_2028_),
    .B2(_2038_),
    .ZN(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2596_ (.I(_2039_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2597_ (.I(\t2pre[7] ),
    .Z(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2598_ (.A1(\t0_top[7] ),
    .A2(_1886_),
    .B1(_1900_),
    .B2(_2040_),
    .ZN(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2599_ (.A1(\t2pre[15] ),
    .A2(_1851_),
    .B1(_1875_),
    .B2(\t2_top[15] ),
    .ZN(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2600_ (.A1(\t1pre[15] ),
    .A2(_1870_),
    .B1(_1842_),
    .B2(\t1_capture[15] ),
    .ZN(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2601_ (.A1(_2041_),
    .A2(_2042_),
    .A3(_2043_),
    .ZN(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2602_ (.A1(\t0pre[7] ),
    .A2(_1919_),
    .B1(_1916_),
    .B2(\t2_capture[7] ),
    .C(_2044_),
    .ZN(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2603_ (.A1(\pw2[7] ),
    .A2(_1880_),
    .B1(_1818_),
    .B2(\t1_capture[7] ),
    .ZN(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2604_ (.A1(\t2_top[7] ),
    .A2(_1994_),
    .B1(_1873_),
    .B2(\t0_capture[7] ),
    .ZN(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2605_ (.A1(\t1_top[15] ),
    .A2(_1902_),
    .B1(_1892_),
    .B2(\t2_capture[15] ),
    .ZN(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2606_ (.A1(_2046_),
    .A2(_2047_),
    .A3(_2048_),
    .ZN(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2607_ (.A1(\t0_top[15] ),
    .A2(_1862_),
    .B1(_1833_),
    .B2(\t0pre[15] ),
    .C(_2049_),
    .ZN(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2608_ (.A1(\t1_top[7] ),
    .A2(_1996_),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2609_ (.A1(\pw1[7] ),
    .A2(_1904_),
    .B1(_1893_),
    .B2(\t1pre[7] ),
    .ZN(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2610_ (.A1(_1867_),
    .A2(_2051_),
    .A3(_2052_),
    .ZN(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2611_ (.A1(\pw0[7] ),
    .A2(_1921_),
    .B1(_1898_),
    .B2(\t0_capture[15] ),
    .C(_2053_),
    .ZN(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2612_ (.A1(_2045_),
    .A2(_2050_),
    .A3(_2054_),
    .ZN(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2613_ (.A1(net27),
    .A2(_1911_),
    .B(_2055_),
    .ZN(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2614_ (.I(_2056_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2615_ (.I(\settings[0] ),
    .ZN(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2616_ (.I(\t0pre[14] ),
    .ZN(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2617_ (.I(\t0pre_counter[12] ),
    .Z(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2618_ (.A1(\t0pre_counter[13] ),
    .A2(_2059_),
    .ZN(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2619_ (.I(\t0pre_counter[2] ),
    .Z(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2620_ (.I(\t0pre_counter[0] ),
    .Z(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2621_ (.A1(\t0pre_counter[3] ),
    .A2(_2061_),
    .A3(\t0pre_counter[1] ),
    .A4(_2062_),
    .ZN(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2622_ (.A1(\t0pre_counter[7] ),
    .A2(\t0pre_counter[6] ),
    .A3(\t0pre_counter[5] ),
    .A4(\t0pre_counter[4] ),
    .ZN(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2623_ (.I(_2064_),
    .Z(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2624_ (.A1(\t0pre_counter[11] ),
    .A2(\t0pre_counter[10] ),
    .A3(\t0pre_counter[9] ),
    .A4(\t0pre_counter[8] ),
    .ZN(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _2625_ (.A1(_2060_),
    .A2(_2063_),
    .A3(_2065_),
    .A4(_2066_),
    .ZN(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2626_ (.A1(\t0pre_counter[14] ),
    .A2(_2067_),
    .Z(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2627_ (.I(\t0pre_counter[14] ),
    .ZN(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2628_ (.I(\t0pre_counter[8] ),
    .Z(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _2629_ (.A1(\t0pre_counter[3] ),
    .A2(\t0pre_counter[2] ),
    .A3(\t0pre_counter[1] ),
    .A4(\t0pre_counter[0] ),
    .Z(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _2630_ (.A1(\t0pre_counter[7] ),
    .A2(\t0pre_counter[6] ),
    .A3(\t0pre_counter[5] ),
    .A4(\t0pre_counter[4] ),
    .Z(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2631_ (.A1(_2070_),
    .A2(_2071_),
    .A3(_2072_),
    .ZN(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2632_ (.I(\t0pre_counter[10] ),
    .Z(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2633_ (.I(\t0pre_counter[9] ),
    .Z(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2634_ (.A1(\t0pre_counter[11] ),
    .A2(_2074_),
    .A3(_2075_),
    .ZN(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2635_ (.A1(_2069_),
    .A2(_2060_),
    .A3(_2073_),
    .A4(_2076_),
    .ZN(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2636_ (.A1(\t0pre_counter[15] ),
    .A2(_2077_),
    .Z(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2637_ (.I(\t0pre[15] ),
    .ZN(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _2638_ (.A1(_2058_),
    .A2(_2068_),
    .B1(_2078_),
    .B2(_2079_),
    .ZN(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _2639_ (.A1(\t0pre_counter[15] ),
    .A2(_2077_),
    .ZN(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2640_ (.I(\t0pre_counter[12] ),
    .ZN(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _2641_ (.A1(_2082_),
    .A2(_2063_),
    .A3(_2064_),
    .A4(_2066_),
    .Z(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2642_ (.A1(\t0pre_counter[13] ),
    .A2(_2083_),
    .ZN(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2643_ (.I(\t0pre[13] ),
    .ZN(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2644_ (.A1(_2058_),
    .A2(_2068_),
    .B1(_2084_),
    .B2(_2085_),
    .ZN(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2645_ (.A1(\t0pre_counter[13] ),
    .A2(_2083_),
    .Z(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2646_ (.A1(_2063_),
    .A2(_2064_),
    .A3(_2066_),
    .ZN(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2647_ (.A1(_2059_),
    .A2(\t0pre[12] ),
    .A3(_2088_),
    .Z(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2648_ (.A1(\t0pre[13] ),
    .A2(_2087_),
    .B(_2089_),
    .ZN(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2649_ (.A1(\t0pre[15] ),
    .A2(_2081_),
    .B(_2086_),
    .C(_2090_),
    .ZN(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2650_ (.I(\t0pre[11] ),
    .ZN(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2651_ (.I(_2088_),
    .Z(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2652_ (.I(_2075_),
    .ZN(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2653_ (.I(_2070_),
    .ZN(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2654_ (.I(_2063_),
    .Z(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _2655_ (.A1(_2094_),
    .A2(_2095_),
    .A3(_2096_),
    .A4(_2065_),
    .ZN(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2656_ (.A1(_2074_),
    .A2(_2097_),
    .B(\t0pre_counter[11] ),
    .ZN(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2657_ (.A1(_2093_),
    .A2(_2098_),
    .ZN(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2658_ (.A1(_2075_),
    .A2(_2070_),
    .A3(_2071_),
    .A4(_2072_),
    .ZN(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2659_ (.A1(_2074_),
    .A2(_2100_),
    .Z(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2660_ (.A1(\t0pre[10] ),
    .A2(_2101_),
    .ZN(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2661_ (.A1(_2092_),
    .A2(_2099_),
    .B(_2102_),
    .ZN(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2662_ (.A1(_2095_),
    .A2(_2096_),
    .A3(_2065_),
    .B(_2094_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2663_ (.A1(_2100_),
    .A2(_0319_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2664_ (.A1(\t0pre[10] ),
    .A2(_2101_),
    .B1(_0320_),
    .B2(\t0pre[9] ),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2665_ (.I(\t0pre[9] ),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2666_ (.A1(_2100_),
    .A2(_0319_),
    .B(_0322_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2667_ (.A1(_2096_),
    .A2(_2065_),
    .B(_2095_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2668_ (.I(\t0pre[8] ),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2669_ (.A1(_2073_),
    .A2(_0324_),
    .B(_0325_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2670_ (.A1(_0323_),
    .A2(_0326_),
    .Z(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2671_ (.A1(_2073_),
    .A2(_0324_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2672_ (.A1(\t0pre[11] ),
    .A2(_2093_),
    .A3(_2098_),
    .B1(_0328_),
    .B2(\t0pre[8] ),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2673_ (.A1(_0321_),
    .A2(_0327_),
    .A3(_0329_),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _2674_ (.A1(_2080_),
    .A2(_2091_),
    .A3(_2103_),
    .A4(_0330_),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2675_ (.I(\t0pre[7] ),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2676_ (.I(_2071_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2677_ (.I(\t0pre_counter[6] ),
    .Z(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2678_ (.I(\t0pre_counter[5] ),
    .Z(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2679_ (.I(\t0pre_counter[4] ),
    .Z(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2680_ (.A1(_0334_),
    .A2(_0335_),
    .A3(_0336_),
    .A4(_0333_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2681_ (.I(\t0pre_counter[7] ),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2682_ (.A1(_0333_),
    .A2(_2072_),
    .B1(_0337_),
    .B2(_0338_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2683_ (.I(_0339_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2684_ (.A1(_0332_),
    .A2(_0340_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2685_ (.A1(_0336_),
    .A2(_0333_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2686_ (.A1(_0335_),
    .A2(_0342_),
    .Z(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2687_ (.A1(_0336_),
    .A2(_2096_),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2688_ (.A1(_2007_),
    .A2(_0343_),
    .B1(_0344_),
    .B2(_1987_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2689_ (.A1(\t0pre_counter[5] ),
    .A2(\t0pre_counter[4] ),
    .A3(_0333_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2690_ (.A1(_0334_),
    .A2(_0346_),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _2691_ (.A1(\t0pre[6] ),
    .A2(_0347_),
    .B1(_0343_),
    .B2(_2007_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _2692_ (.A1(_0334_),
    .A2(_0346_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2693_ (.I(\t0pre[6] ),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _2694_ (.A1(_0332_),
    .A2(_0340_),
    .B1(_0345_),
    .B2(_0348_),
    .C1(_0349_),
    .C2(_0350_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2695_ (.A1(_0332_),
    .A2(_0339_),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2696_ (.A1(_0332_),
    .A2(_0340_),
    .B1(_0349_),
    .B2(_0350_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2697_ (.I(\t0pre[5] ),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2698_ (.A1(_0335_),
    .A2(_0342_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2699_ (.A1(_1987_),
    .A2(_0344_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2700_ (.A1(\t0pre[4] ),
    .A2(_0344_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2701_ (.A1(_0354_),
    .A2(_0355_),
    .B(_0356_),
    .C(_0357_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2702_ (.A1(_0352_),
    .A2(_0353_),
    .A3(_0348_),
    .A4(_0358_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2703_ (.I(\t0pre_counter[1] ),
    .Z(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2704_ (.A1(_2061_),
    .A2(_0360_),
    .A3(_2062_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2705_ (.A1(\t0pre_counter[3] ),
    .A2(_0361_),
    .Z(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2706_ (.I(_2062_),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2707_ (.A1(_0360_),
    .A2(_0363_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2708_ (.A1(_2061_),
    .A2(_0364_),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2709_ (.A1(\t0pre[3] ),
    .A2(_0362_),
    .B1(_0365_),
    .B2(_1945_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2710_ (.A1(_0360_),
    .A2(_2062_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2711_ (.A1(\t0pre[1] ),
    .A2(_0367_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2712_ (.A1(\t0pre[1] ),
    .A2(_0367_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2713_ (.A1(_0363_),
    .A2(\t0pre[0] ),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2714_ (.A1(_0368_),
    .A2(_0369_),
    .A3(_0370_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2715_ (.A1(_1945_),
    .A2(_0365_),
    .B1(_0368_),
    .B2(_0371_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2716_ (.A1(\t0pre[3] ),
    .A2(_0362_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2717_ (.A1(_0366_),
    .A2(_0372_),
    .B(_0373_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2718_ (.A1(_0341_),
    .A2(_0351_),
    .B1(_0359_),
    .B2(_0374_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2719_ (.A1(_0323_),
    .A2(_0326_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2720_ (.A1(_0321_),
    .A2(_0376_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2721_ (.A1(\t0pre[11] ),
    .A2(_2093_),
    .A3(_2098_),
    .B1(_2103_),
    .B2(_0377_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2722_ (.A1(_2080_),
    .A2(_2091_),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2723_ (.A1(_2059_),
    .A2(_2093_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2724_ (.I(\t0pre[12] ),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2725_ (.A1(_2085_),
    .A2(_2084_),
    .B1(_0380_),
    .B2(_0381_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2726_ (.A1(_2086_),
    .A2(_0382_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2727_ (.A1(\t0pre[15] ),
    .A2(_2081_),
    .B1(_2080_),
    .B2(_0383_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _2728_ (.A1(_0331_),
    .A2(_0375_),
    .B1(_0378_),
    .B2(_0379_),
    .C(_0384_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2729_ (.A1(_2080_),
    .A2(_2091_),
    .A3(_2103_),
    .A4(_0330_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2730_ (.I(_0365_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2731_ (.I(\t0pre[2] ),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2732_ (.A1(_0363_),
    .A2(\t0pre[0] ),
    .B1(_0387_),
    .B2(_0388_),
    .C(_0373_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2733_ (.A1(_0359_),
    .A2(_0366_),
    .A3(_0371_),
    .A4(_0389_),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2734_ (.A1(\t0pre_counter[15] ),
    .A2(_2077_),
    .B1(_0386_),
    .B2(_0390_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2735_ (.I(last_tmr0_clk),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2736_ (.I(tmr0_ext),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2737_ (.A1(net18),
    .A2(_0392_),
    .B(_0393_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2738_ (.A1(_0385_),
    .A2(_0391_),
    .B(_0394_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2739_ (.I(_0395_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2740_ (.I(\t0_top[7] ),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2741_ (.I(\timer0[7] ),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2742_ (.I(\timer0[6] ),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2743_ (.I(\t0_top[6] ),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _2744_ (.I(\timer0[6] ),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _2745_ (.I(\timer0[5] ),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2746_ (.I(\t0_top[5] ),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2747_ (.I(\t0_top[4] ),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2748_ (.I(\timer0[4] ),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2749_ (.I(\timer0[3] ),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2750_ (.I(\t0_top[2] ),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2751_ (.I(\timer0[1] ),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2752_ (.I(\timer0[0] ),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2753_ (.A1(\t0_top[1] ),
    .A2(_0408_),
    .B(_0409_),
    .C(\t0_top[0] ),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2754_ (.I(\timer0[2] ),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2755_ (.A1(\t0_top[2] ),
    .A2(_0411_),
    .B1(_0408_),
    .B2(\t0_top[1] ),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2756_ (.A1(\t0_top[3] ),
    .A2(_0406_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2757_ (.A1(_0407_),
    .A2(\timer0[2] ),
    .B1(_0410_),
    .B2(_0412_),
    .C(_0413_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2758_ (.A1(\t0_top[4] ),
    .A2(_0405_),
    .B1(_0406_),
    .B2(\t0_top[3] ),
    .C(_0414_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2759_ (.A1(_0403_),
    .A2(\timer0[5] ),
    .B1(\timer0[4] ),
    .B2(_0404_),
    .C(_0415_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2760_ (.A1(\t0_top[6] ),
    .A2(_0401_),
    .B1(_0402_),
    .B2(\t0_top[5] ),
    .C(_0416_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2761_ (.A1(_0397_),
    .A2(_0398_),
    .B1(_0399_),
    .B2(_0400_),
    .C(_0417_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2762_ (.I(\t0_top[11] ),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2763_ (.I(\timer0[10] ),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2764_ (.I(\t0_top[10] ),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2765_ (.A1(_0419_),
    .A2(\timer0[11] ),
    .B1(_0420_),
    .B2(_0421_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2766_ (.I(\timer0[9] ),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2767_ (.I(\timer0[8] ),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2768_ (.A1(\t0_top[9] ),
    .A2(_0423_),
    .B1(_0424_),
    .B2(\t0_top[8] ),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2769_ (.I(_0425_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2770_ (.I(\timer0[10] ),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2771_ (.A1(\t0_top[10] ),
    .A2(_0427_),
    .B1(_0423_),
    .B2(\t0_top[9] ),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2772_ (.A1(_0422_),
    .A2(_0426_),
    .A3(_0428_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2773_ (.I(\t0_top[8] ),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2774_ (.I(\timer0[14] ),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2775_ (.A1(\t0_top[14] ),
    .A2(_0431_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2776_ (.A1(_0430_),
    .A2(\timer0[8] ),
    .B1(\timer0[7] ),
    .B2(_0397_),
    .C(_0432_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2777_ (.I(\timer0[15] ),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2778_ (.A1(\t0_top[15] ),
    .A2(_0434_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2779_ (.I(\timer0[13] ),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2780_ (.A1(\t0_top[13] ),
    .A2(_0436_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2781_ (.I(\t0_top[15] ),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2782_ (.I(\timer0[14] ),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2783_ (.I(\t0_top[14] ),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2784_ (.A1(_0438_),
    .A2(\timer0[15] ),
    .B1(_0439_),
    .B2(_0440_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2785_ (.I(\timer0[12] ),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2786_ (.A1(\t0_top[13] ),
    .A2(_0436_),
    .B1(_0442_),
    .B2(\t0_top[12] ),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2787_ (.I(\t0_top[12] ),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2788_ (.A1(_0444_),
    .A2(\timer0[12] ),
    .B1(\timer0[11] ),
    .B2(_0419_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2789_ (.A1(_0443_),
    .A2(_0445_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2790_ (.A1(_0435_),
    .A2(_0437_),
    .A3(_0441_),
    .A4(_0446_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2791_ (.A1(_0429_),
    .A2(_0433_),
    .A3(_0447_),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2792_ (.A1(_0425_),
    .A2(_0428_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2793_ (.A1(_0422_),
    .A2(_0449_),
    .B(_0445_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2794_ (.A1(_0443_),
    .A2(_0450_),
    .B(_0432_),
    .C(_0437_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2795_ (.A1(_0451_),
    .A2(_0441_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2796_ (.A1(_0435_),
    .A2(_0452_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _2797_ (.A1(_0418_),
    .A2(_0448_),
    .B(_0453_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2798_ (.A1(_0396_),
    .A2(_0454_),
    .Z(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2799_ (.I(_0455_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2800_ (.I(net12),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2801_ (.A1(net8),
    .A2(net7),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2802_ (.I(_0458_),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2803_ (.I(_0459_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2804_ (.A1(_1822_),
    .A2(_1844_),
    .A3(_0460_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2805_ (.A1(_0457_),
    .A2(_0461_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2806_ (.I(_1802_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2807_ (.I(_0463_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2808_ (.I(_0464_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2809_ (.A1(net28),
    .A2(_0456_),
    .B(_0462_),
    .C(_0465_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2810_ (.A1(_2057_),
    .A2(_0456_),
    .B(_0466_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2811_ (.I(_1803_),
    .Z(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2812_ (.I(_0467_),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2813_ (.I(net13),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2814_ (.A1(_0469_),
    .A2(_0461_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2815_ (.I(last_tmr1_clk),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2816_ (.I(tmr1_ext),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2817_ (.A1(net19),
    .A2(_0471_),
    .B(_0472_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2818_ (.I(\t1pre_counter[14] ),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2819_ (.A1(\t1pre_counter[13] ),
    .A2(\t1pre_counter[12] ),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2820_ (.I(\t1pre_counter[2] ),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2821_ (.A1(\t1pre_counter[3] ),
    .A2(_0476_),
    .A3(\t1pre_counter[1] ),
    .A4(\t1pre_counter[0] ),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2822_ (.A1(\t1pre_counter[7] ),
    .A2(\t1pre_counter[6] ),
    .A3(\t1pre_counter[5] ),
    .A4(\t1pre_counter[4] ),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2823_ (.A1(\t1pre_counter[11] ),
    .A2(\t1pre_counter[10] ),
    .A3(\t1pre_counter[9] ),
    .A4(\t1pre_counter[8] ),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2824_ (.A1(_0475_),
    .A2(_0477_),
    .A3(_0478_),
    .A4(_0479_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2825_ (.A1(_0474_),
    .A2(_0480_),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2826_ (.A1(\t1pre_counter[14] ),
    .A2(_0480_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2827_ (.A1(\t1pre_counter[15] ),
    .A2(_0482_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2828_ (.A1(\t1pre[14] ),
    .A2(_0481_),
    .B1(_0483_),
    .B2(\t1pre[15] ),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2829_ (.I(\t1pre[15] ),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2830_ (.A1(\t1pre_counter[15] ),
    .A2(_0482_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2831_ (.I(\t1pre_counter[12] ),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2832_ (.A1(_0487_),
    .A2(_0477_),
    .A3(_0478_),
    .A4(_0479_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2833_ (.A1(\t1pre_counter[13] ),
    .A2(_0488_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2834_ (.A1(\t1pre[14] ),
    .A2(_0481_),
    .B1(_0489_),
    .B2(\t1pre[13] ),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2835_ (.I(\t1pre[13] ),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2836_ (.A1(\t1pre_counter[13] ),
    .A2(_0488_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2837_ (.A1(_0477_),
    .A2(_0478_),
    .A3(_0479_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2838_ (.A1(_0487_),
    .A2(\t1pre[12] ),
    .A3(_0493_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2839_ (.A1(_0491_),
    .A2(_0492_),
    .B(_0494_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2840_ (.A1(_0485_),
    .A2(_0486_),
    .B(_0490_),
    .C(_0495_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2841_ (.I(\t1pre_counter[10] ),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2842_ (.I(\t1pre_counter[8] ),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2843_ (.A1(\t1pre_counter[3] ),
    .A2(\t1pre_counter[2] ),
    .A3(\t1pre_counter[1] ),
    .A4(\t1pre_counter[0] ),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2844_ (.A1(\t1pre_counter[7] ),
    .A2(\t1pre_counter[6] ),
    .A3(\t1pre_counter[5] ),
    .A4(\t1pre_counter[4] ),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2845_ (.A1(\t1pre_counter[9] ),
    .A2(_0498_),
    .A3(_0499_),
    .A4(_0500_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2846_ (.A1(_0497_),
    .A2(_0501_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2847_ (.A1(\t1pre[10] ),
    .A2(_0502_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2848_ (.I(_0493_),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2849_ (.A1(_0497_),
    .A2(_0501_),
    .B(\t1pre_counter[11] ),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2850_ (.A1(_0504_),
    .A2(_0505_),
    .B(_1972_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2851_ (.A1(_0503_),
    .A2(_0506_),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2852_ (.I(\t1pre_counter[9] ),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2853_ (.A1(\t1pre_counter[8] ),
    .A2(_0499_),
    .A3(_0500_),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2854_ (.A1(_0508_),
    .A2(_0509_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2855_ (.A1(\t1pre[10] ),
    .A2(_0502_),
    .B1(_0510_),
    .B2(_1929_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2856_ (.I(\t1pre[9] ),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2857_ (.A1(_0508_),
    .A2(_0509_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2858_ (.I(_0499_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2859_ (.A1(_0514_),
    .A2(_0500_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2860_ (.A1(_0498_),
    .A2(_0515_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2861_ (.I(\t1pre[8] ),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2862_ (.A1(_0512_),
    .A2(_0513_),
    .B1(_0516_),
    .B2(_0517_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2863_ (.A1(_0498_),
    .A2(_0515_),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2864_ (.A1(\t1pre[11] ),
    .A2(_0504_),
    .A3(_0505_),
    .B1(_0519_),
    .B2(\t1pre[8] ),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2865_ (.A1(_0511_),
    .A2(_0518_),
    .A3(_0520_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2866_ (.A1(_0484_),
    .A2(_0496_),
    .A3(_0507_),
    .A4(_0521_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2867_ (.I(\t1pre_counter[6] ),
    .Z(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2868_ (.I(\t1pre_counter[5] ),
    .Z(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2869_ (.I(\t1pre_counter[4] ),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2870_ (.A1(_0523_),
    .A2(_0524_),
    .A3(_0525_),
    .A4(_0514_),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2871_ (.A1(\t1pre_counter[7] ),
    .A2(_0526_),
    .B(_0515_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2872_ (.A1(\t1pre[7] ),
    .A2(_0527_),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2873_ (.A1(_0525_),
    .A2(_0514_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2874_ (.A1(_0524_),
    .A2(_0529_),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2875_ (.A1(_0525_),
    .A2(_0477_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2876_ (.A1(\t1pre[4] ),
    .A2(_0531_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2877_ (.A1(_2012_),
    .A2(_0530_),
    .B(_0532_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2878_ (.A1(\t1pre_counter[5] ),
    .A2(\t1pre_counter[4] ),
    .A3(_0514_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2879_ (.A1(_0523_),
    .A2(_0534_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2880_ (.A1(_2030_),
    .A2(_0535_),
    .B1(_0530_),
    .B2(_2012_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2881_ (.A1(\t1pre[7] ),
    .A2(_0527_),
    .B1(_0535_),
    .B2(_2030_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2882_ (.A1(_0533_),
    .A2(_0536_),
    .B(_0537_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2883_ (.I(\t1pre[6] ),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2884_ (.A1(_0523_),
    .A2(_0534_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2885_ (.A1(_0524_),
    .A2(_0529_),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2886_ (.I(\t1pre[5] ),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2887_ (.A1(_0539_),
    .A2(_0540_),
    .B1(_0541_),
    .B2(_0542_),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2888_ (.A1(\t1pre[4] ),
    .A2(_0531_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2889_ (.A1(\t1pre[5] ),
    .A2(_0530_),
    .B(_0532_),
    .C(_0544_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2890_ (.A1(_0528_),
    .A2(_0537_),
    .A3(_0543_),
    .A4(_0545_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2891_ (.I(\t1pre_counter[1] ),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2892_ (.I(\t1pre_counter[0] ),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2893_ (.A1(_0476_),
    .A2(_0547_),
    .A3(_0548_),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2894_ (.A1(\t1pre_counter[3] ),
    .A2(_0549_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2895_ (.A1(_0547_),
    .A2(_0548_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2896_ (.A1(_0476_),
    .A2(_0551_),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2897_ (.A1(\t1pre[3] ),
    .A2(_0550_),
    .B1(_0552_),
    .B2(_1951_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2898_ (.A1(_0547_),
    .A2(_0548_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2899_ (.A1(\t1pre[1] ),
    .A2(_0554_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2900_ (.I(_0548_),
    .Z(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2901_ (.A1(_0556_),
    .A2(\t1pre[0] ),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2902_ (.A1(\t1pre[1] ),
    .A2(_0554_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2903_ (.A1(_0555_),
    .A2(_0557_),
    .B(_0558_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2904_ (.A1(_1951_),
    .A2(_0552_),
    .B(_0559_),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2905_ (.A1(\t1pre[3] ),
    .A2(_0550_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2906_ (.A1(_0553_),
    .A2(_0560_),
    .B(_0561_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2907_ (.A1(_0528_),
    .A2(_0538_),
    .B1(_0546_),
    .B2(_0562_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2908_ (.A1(_0487_),
    .A2(_0504_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2909_ (.A1(\t1pre[13] ),
    .A2(_0489_),
    .B1(_0564_),
    .B2(\t1pre[12] ),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2910_ (.A1(_0490_),
    .A2(_0565_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2911_ (.A1(_0484_),
    .A2(_0566_),
    .Z(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2912_ (.A1(\t1pre[15] ),
    .A2(_0483_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2913_ (.A1(_0504_),
    .A2(_0505_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2914_ (.A1(_1972_),
    .A2(_0569_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2915_ (.A1(_1929_),
    .A2(_0510_),
    .B1(_0519_),
    .B2(\t1pre[8] ),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2916_ (.A1(_0511_),
    .A2(_0571_),
    .B(_0503_),
    .C(_0506_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2917_ (.A1(_0484_),
    .A2(_0496_),
    .A3(_0570_),
    .A4(_0572_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _2918_ (.A1(_0522_),
    .A2(_0563_),
    .B1(_0567_),
    .B2(_0568_),
    .C(_0573_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2919_ (.A1(\t1pre_counter[11] ),
    .A2(_0497_),
    .A3(_0508_),
    .A4(_0509_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2920_ (.A1(_0474_),
    .A2(_0475_),
    .A3(_0575_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2921_ (.A1(_0484_),
    .A2(_0496_),
    .A3(_0507_),
    .A4(_0521_),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2922_ (.A1(_0556_),
    .A2(_1895_),
    .B(_0558_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2923_ (.A1(_0556_),
    .A2(_1895_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2924_ (.A1(\t1pre[2] ),
    .A2(_0552_),
    .B(_0579_),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2925_ (.A1(_0561_),
    .A2(_0555_),
    .A3(_0578_),
    .A4(_0580_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2926_ (.A1(_0546_),
    .A2(_0553_),
    .A3(_0581_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2927_ (.A1(\t1pre_counter[15] ),
    .A2(_0576_),
    .B1(_0577_),
    .B2(_0582_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _2928_ (.A1(_0574_),
    .A2(_0583_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2929_ (.I(\timer1[15] ),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2930_ (.A1(\t1_top[15] ),
    .A2(_0585_),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2931_ (.I(\t1_top[14] ),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2932_ (.I(\timer1[14] ),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2933_ (.I(\timer1[13] ),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2934_ (.A1(\t1_top[13] ),
    .A2(_0589_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2935_ (.I(\t1_top[12] ),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2936_ (.I(\timer1[12] ),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2937_ (.I(\t1_top[11] ),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2938_ (.A1(_0591_),
    .A2(_0592_),
    .B1(\timer1[11] ),
    .B2(_0593_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2939_ (.I(\timer1[9] ),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2940_ (.I(_0595_),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2941_ (.I(\timer1[8] ),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2942_ (.A1(\t1_top[9] ),
    .A2(_0596_),
    .B1(_0597_),
    .B2(\t1_top[8] ),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2943_ (.I(\timer1[10] ),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2944_ (.I(_0599_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2945_ (.A1(\t1_top[10] ),
    .A2(_0600_),
    .B1(_0595_),
    .B2(\t1_top[9] ),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2946_ (.I(\timer1[11] ),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2947_ (.A1(\t1_top[11] ),
    .A2(_0602_),
    .B1(_0599_),
    .B2(\t1_top[10] ),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2948_ (.A1(_0598_),
    .A2(_0601_),
    .B(_0603_),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2949_ (.I(\t1_top[13] ),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2950_ (.A1(_0605_),
    .A2(\timer1[13] ),
    .B1(\timer1[12] ),
    .B2(_0591_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2951_ (.A1(_0594_),
    .A2(_0604_),
    .B(_0606_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2952_ (.A1(_0587_),
    .A2(_0588_),
    .B(_0590_),
    .C(_0607_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2953_ (.I(\t1_top[15] ),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2954_ (.A1(_0609_),
    .A2(\timer1[15] ),
    .B1(\timer1[14] ),
    .B2(_0587_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2955_ (.A1(_0608_),
    .A2(_0610_),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2956_ (.I(\timer1[6] ),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2957_ (.I(\t1_top[4] ),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2958_ (.I(\timer1[2] ),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _2959_ (.I(\timer1[1] ),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2960_ (.I(\t1_top[1] ),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2961_ (.I(\timer1[1] ),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2962_ (.I(\t1_top[0] ),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2963_ (.A1(_0616_),
    .A2(_0617_),
    .B(\timer1[0] ),
    .C(_0618_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2964_ (.A1(\t1_top[2] ),
    .A2(_0614_),
    .B1(_0615_),
    .B2(\t1_top[1] ),
    .C(_0619_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2965_ (.I(\timer1[3] ),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2966_ (.A1(\t1_top[3] ),
    .A2(_0621_),
    .B1(_0614_),
    .B2(\t1_top[2] ),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2967_ (.A1(\t1_top[3] ),
    .A2(_0621_),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2968_ (.A1(_0613_),
    .A2(\timer1[4] ),
    .B1(_0620_),
    .B2(_0622_),
    .C(_0623_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2969_ (.I(\t1_top[5] ),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2970_ (.I(\timer1[4] ),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2971_ (.A1(_0625_),
    .A2(\timer1[5] ),
    .B1(_0626_),
    .B2(_0613_),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2972_ (.I(\timer1[5] ),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2973_ (.A1(\t1_top[6] ),
    .A2(_0612_),
    .B1(_0624_),
    .B2(_0627_),
    .C1(_0628_),
    .C2(\t1_top[5] ),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2974_ (.I(\timer1[7] ),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2975_ (.I(_0630_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2976_ (.A1(\t1_top[7] ),
    .A2(_0631_),
    .B1(_0612_),
    .B2(\t1_top[6] ),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2977_ (.A1(_0629_),
    .A2(_0632_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2978_ (.A1(_0603_),
    .A2(_0598_),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2979_ (.I(_0588_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2980_ (.A1(\t1_top[14] ),
    .A2(_0635_),
    .B1(_0597_),
    .B2(\t1_top[8] ),
    .C1(_0630_),
    .C2(\t1_top[7] ),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2981_ (.I(_0606_),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2982_ (.A1(_0586_),
    .A2(_0590_),
    .A3(_0610_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2983_ (.A1(_0637_),
    .A2(_0594_),
    .A3(_0638_),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2984_ (.A1(_0601_),
    .A2(_0634_),
    .A3(_0636_),
    .A4(_0639_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2985_ (.A1(_0586_),
    .A2(_0611_),
    .B1(_0633_),
    .B2(_0640_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _2986_ (.A1(_0473_),
    .A2(_0584_),
    .A3(_0641_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2987_ (.I0(\settings[1] ),
    .I1(net29),
    .S(_0642_),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2988_ (.A1(_0468_),
    .A2(_0470_),
    .A3(_0643_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2989_ (.I(_0644_),
    .Z(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2990_ (.A1(net34),
    .A2(_0456_),
    .B(_1805_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2991_ (.A1(net34),
    .A2(_0456_),
    .B(_0645_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2992_ (.I(_0467_),
    .Z(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2993_ (.A1(net35),
    .A2(_0642_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2994_ (.A1(_0646_),
    .A2(_0647_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2995_ (.I(_0648_),
    .Z(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2996_ (.I(\pwm_ctr0[5] ),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2997_ (.A1(\pw0[5] ),
    .A2(_0649_),
    .B(_0465_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2998_ (.I(\pw0[4] ),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2999_ (.I(\pwm_ctr0[6] ),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3000_ (.I(\pw0[6] ),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3001_ (.I(\pwm_ctr0[0] ),
    .Z(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3002_ (.A1(\pw0[0] ),
    .A2(_0654_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _3003_ (.A1(_0651_),
    .A2(\pwm_ctr0[4] ),
    .B1(_0652_),
    .B2(_0653_),
    .C(_0655_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3004_ (.I(\pwm_ctr0[3] ),
    .Z(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3005_ (.I(_0657_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3006_ (.I(\pwm_ctr0[7] ),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3007_ (.A1(\pw0[3] ),
    .A2(_0658_),
    .B1(\pwm_ctr0[4] ),
    .B2(_0651_),
    .C1(\pw0[7] ),
    .C2(_0659_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3008_ (.I(\pw0[7] ),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3009_ (.I(\pw0[2] ),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3010_ (.A1(_0662_),
    .A2(\pwm_ctr0[2] ),
    .B1(_0658_),
    .B2(\pw0[3] ),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3011_ (.A1(\pw0[5] ),
    .A2(_0649_),
    .B1(\pwm_ctr0[7] ),
    .B2(_0661_),
    .C(_0663_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3012_ (.A1(\pw0[1] ),
    .A2(\pwm_ctr0[1] ),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3013_ (.A1(_0662_),
    .A2(\pwm_ctr0[2] ),
    .B1(\pwm_ctr0[6] ),
    .B2(_0653_),
    .C(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3014_ (.A1(_0660_),
    .A2(_0664_),
    .A3(_0666_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3015_ (.A1(\pwm_ctr0[0] ),
    .A2(\pwm_ctr0[1] ),
    .A3(\pwm_ctr0[2] ),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3016_ (.A1(\pwm_ctr0[3] ),
    .A2(\pwm_ctr0[4] ),
    .A3(_0668_),
    .Z(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3017_ (.A1(\pwm_ctr0[5] ),
    .A2(_0669_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3018_ (.A1(_0652_),
    .A2(\pwm_ctr0[7] ),
    .A3(_0670_),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3019_ (.A1(_1781_),
    .A2(_0671_),
    .B(net31),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3020_ (.A1(_0650_),
    .A2(_0656_),
    .A3(_0667_),
    .B(_0672_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3021_ (.I(\pwm_ctr1[5] ),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3022_ (.A1(\pw1[5] ),
    .A2(_0673_),
    .B(_0467_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3023_ (.I(\pw1[4] ),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3024_ (.I(\pwm_ctr1[6] ),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3025_ (.I(\pw1[6] ),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3026_ (.I(\pwm_ctr1[0] ),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3027_ (.A1(\pw1[0] ),
    .A2(_0678_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _3028_ (.A1(_0675_),
    .A2(\pwm_ctr1[4] ),
    .B1(_0676_),
    .B2(_0677_),
    .C(_0679_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3029_ (.I(\pwm_ctr1[3] ),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3030_ (.I(_0681_),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3031_ (.I(\pwm_ctr1[7] ),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3032_ (.A1(\pw1[3] ),
    .A2(_0682_),
    .B1(\pwm_ctr1[4] ),
    .B2(_0675_),
    .C1(\pw1[7] ),
    .C2(_0683_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3033_ (.I(\pw1[7] ),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3034_ (.I(\pw1[2] ),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3035_ (.A1(_0686_),
    .A2(\pwm_ctr1[2] ),
    .B1(_0682_),
    .B2(\pw1[3] ),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3036_ (.A1(\pw1[5] ),
    .A2(_0673_),
    .B1(\pwm_ctr1[7] ),
    .B2(_0685_),
    .C(_0687_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3037_ (.A1(\pw1[1] ),
    .A2(\pwm_ctr1[1] ),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3038_ (.A1(_0686_),
    .A2(\pwm_ctr1[2] ),
    .B1(\pwm_ctr1[6] ),
    .B2(_0677_),
    .C(_0689_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3039_ (.A1(_0684_),
    .A2(_0688_),
    .A3(_0690_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3040_ (.A1(\pwm_ctr1[0] ),
    .A2(\pwm_ctr1[1] ),
    .A3(\pwm_ctr1[2] ),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3041_ (.A1(\pwm_ctr1[3] ),
    .A2(\pwm_ctr1[4] ),
    .A3(_0692_),
    .Z(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3042_ (.A1(\pwm_ctr1[5] ),
    .A2(_0693_),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3043_ (.A1(_0676_),
    .A2(\pwm_ctr1[7] ),
    .A3(_0694_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3044_ (.A1(_1781_),
    .A2(_0695_),
    .B(net32),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3045_ (.A1(_0674_),
    .A2(_0680_),
    .A3(_0691_),
    .B(_0696_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3046_ (.I(\pw2[0] ),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3047_ (.I(\pw2[6] ),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3048_ (.A1(_0697_),
    .A2(_1778_),
    .B1(_1786_),
    .B2(\pw2[1] ),
    .C1(_0698_),
    .C2(\pwm_ctr2[6] ),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3049_ (.I(\pw2[2] ),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3050_ (.A1(_0700_),
    .A2(\pwm_ctr2[2] ),
    .B1(\pwm_ctr2[6] ),
    .B2(_0698_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3051_ (.I(\pw2[4] ),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3052_ (.A1(\pw2[1] ),
    .A2(_1786_),
    .B1(\pwm_ctr2[4] ),
    .B2(_0702_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3053_ (.A1(_0700_),
    .A2(\pwm_ctr2[2] ),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3054_ (.A1(_0697_),
    .A2(\pwm_ctr2[0] ),
    .B(_0704_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3055_ (.I(\pw2[3] ),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3056_ (.I(\pw2[7] ),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3057_ (.A1(_0706_),
    .A2(\pwm_ctr2[3] ),
    .B1(\pwm_ctr2[7] ),
    .B2(_0707_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _3058_ (.A1(_0701_),
    .A2(_0703_),
    .A3(_0705_),
    .A4(_0708_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3059_ (.A1(_0699_),
    .A2(_0709_),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3060_ (.I(\pwm_ctr2[5] ),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3061_ (.A1(\pw2[5] ),
    .A2(_0711_),
    .B(_1780_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3062_ (.A1(_0706_),
    .A2(\pwm_ctr2[3] ),
    .B1(\pwm_ctr2[4] ),
    .B2(_0702_),
    .C1(_0707_),
    .C2(_1801_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3063_ (.A1(\pw2[5] ),
    .A2(_0711_),
    .B(_0712_),
    .C(_0713_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3064_ (.A1(_1801_),
    .A2(_0465_),
    .A3(_1800_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3065_ (.A1(net33),
    .A2(_0715_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3066_ (.A1(_0710_),
    .A2(_0714_),
    .B(_0716_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3067_ (.I(net14),
    .Z(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3068_ (.A1(net8),
    .A2(net7),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3069_ (.I(_0718_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3070_ (.A1(_1836_),
    .A2(_0719_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _3071_ (.A1(_0717_),
    .A2(net13),
    .A3(net12),
    .A4(_0720_),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3072_ (.A1(\settings[0] ),
    .A2(_0721_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3073_ (.I(net9),
    .Z(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3074_ (.I(_0723_),
    .Z(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3075_ (.A1(net14),
    .A2(net13),
    .A3(net12),
    .A4(_0720_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3076_ (.I(_0725_),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3077_ (.A1(_0724_),
    .A2(_0726_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3078_ (.A1(_0722_),
    .A2(_0727_),
    .B(_1782_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3079_ (.I(net10),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3080_ (.I(_0728_),
    .Z(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3081_ (.A1(\settings[1] ),
    .A2(_0725_),
    .B(_1805_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3082_ (.A1(_0729_),
    .A2(_0726_),
    .B(_0730_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3083_ (.I(net11),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3084_ (.I(_0731_),
    .Z(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3085_ (.I(_1804_),
    .Z(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3086_ (.A1(\settings[2] ),
    .A2(_0725_),
    .B(_0733_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3087_ (.A1(_0732_),
    .A2(_0726_),
    .B(_0734_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3088_ (.I(net15),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3089_ (.I(_0735_),
    .Z(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3090_ (.A1(tmr0_ext),
    .A2(_0725_),
    .B(_0733_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3091_ (.A1(_0736_),
    .A2(_0726_),
    .B(_0737_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3092_ (.I(net16),
    .Z(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3093_ (.A1(_0738_),
    .A2(_0721_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3094_ (.I(_1788_),
    .Z(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3095_ (.A1(_0472_),
    .A2(_0721_),
    .B(_0739_),
    .C(_0740_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3096_ (.I(net30),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3097_ (.I(\t2pre_counter[13] ),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3098_ (.I(\t2pre_counter[12] ),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3099_ (.A1(_0742_),
    .A2(_0743_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3100_ (.A1(\t2pre_counter[3] ),
    .A2(\t2pre_counter[2] ),
    .A3(\t2pre_counter[1] ),
    .A4(\t2pre_counter[0] ),
    .Z(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3101_ (.A1(\t2pre_counter[6] ),
    .A2(\t2pre_counter[5] ),
    .A3(\t2pre_counter[4] ),
    .Z(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3102_ (.A1(\t2pre_counter[11] ),
    .A2(\t2pre_counter[10] ),
    .A3(\t2pre_counter[9] ),
    .A4(\t2pre_counter[8] ),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3103_ (.A1(\t2pre_counter[7] ),
    .A2(_0745_),
    .A3(_0746_),
    .A4(_0747_),
    .Z(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3104_ (.I(_0748_),
    .Z(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3105_ (.A1(_0744_),
    .A2(_0749_),
    .B(\t2pre_counter[14] ),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3106_ (.I(\t2pre_counter[14] ),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3107_ (.A1(\t2pre_counter[13] ),
    .A2(\t2pre_counter[12] ),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3108_ (.I(_0745_),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3109_ (.I(_0746_),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3110_ (.A1(\t2pre_counter[7] ),
    .A2(_0753_),
    .A3(_0754_),
    .A4(_0747_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3111_ (.I(_0755_),
    .Z(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3112_ (.A1(_0751_),
    .A2(_0752_),
    .A3(_0756_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3113_ (.A1(_0750_),
    .A2(_0757_),
    .Z(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3114_ (.I(\t2pre_counter[15] ),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3115_ (.A1(_0751_),
    .A2(_0752_),
    .A3(_0755_),
    .B(_0759_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3116_ (.A1(\t2pre_counter[15] ),
    .A2(\t2pre_counter[14] ),
    .A3(_0744_),
    .A4(_0749_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3117_ (.A1(_0760_),
    .A2(_0761_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3118_ (.A1(\t2pre[14] ),
    .A2(_0758_),
    .B1(_0762_),
    .B2(\t2pre[15] ),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3119_ (.A1(\t2pre_counter[12] ),
    .A2(_0749_),
    .B(\t2pre_counter[13] ),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3120_ (.A1(_0752_),
    .A2(_0755_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_4 _3121_ (.A1(\t2pre[14] ),
    .A2(_0750_),
    .A3(_0757_),
    .B1(_0764_),
    .B2(_0765_),
    .B3(\t2pre[13] ),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3122_ (.I(\t2pre[15] ),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3123_ (.A1(_0767_),
    .A2(_0760_),
    .A3(_0761_),
    .Z(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3124_ (.A1(_0744_),
    .A2(_0749_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3125_ (.A1(_0743_),
    .A2(_0756_),
    .B(_0742_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3126_ (.I(\t2pre[13] ),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3127_ (.A1(_0769_),
    .A2(_0770_),
    .B(_0771_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3128_ (.A1(\t2pre_counter[12] ),
    .A2(_0748_),
    .Z(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3129_ (.A1(\t2pre[12] ),
    .A2(_0773_),
    .Z(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3130_ (.A1(_0766_),
    .A2(_0768_),
    .A3(_0772_),
    .A4(_0774_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3131_ (.I(\t2pre_counter[10] ),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3132_ (.I(\t2pre_counter[9] ),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3133_ (.I(\t2pre_counter[8] ),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3134_ (.I(\t2pre_counter[7] ),
    .Z(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3135_ (.I(_0753_),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3136_ (.I(_0754_),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3137_ (.A1(_0778_),
    .A2(_0779_),
    .A3(_0780_),
    .A4(_0781_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3138_ (.A1(_0776_),
    .A2(_0777_),
    .A3(_0782_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3139_ (.A1(_0778_),
    .A2(_0779_),
    .A3(_0753_),
    .A4(_0754_),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3140_ (.A1(\t2pre_counter[9] ),
    .A2(_0784_),
    .B(\t2pre_counter[10] ),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _3141_ (.A1(_0783_),
    .A2(_0785_),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3142_ (.I(\t2pre_counter[11] ),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3143_ (.A1(_0776_),
    .A2(_0777_),
    .A3(_0782_),
    .B(_0787_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3144_ (.A1(_0756_),
    .A2(_0788_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3145_ (.A1(_1947_),
    .A2(_0786_),
    .B1(_0789_),
    .B2(\t2pre[11] ),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3146_ (.I(\t2pre[11] ),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3147_ (.A1(_0791_),
    .A2(_0756_),
    .A3(_0788_),
    .Z(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3148_ (.A1(_0777_),
    .A2(_0784_),
    .Z(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3149_ (.A1(\t2pre[10] ),
    .A2(_0783_),
    .A3(_0785_),
    .B1(_0793_),
    .B2(_1923_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3150_ (.I(\t2pre[9] ),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3151_ (.A1(\t2pre_counter[9] ),
    .A2(_0784_),
    .Z(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3152_ (.A1(_0779_),
    .A2(_0753_),
    .A3(_0754_),
    .Z(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3153_ (.A1(_0778_),
    .A2(_0797_),
    .Z(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3154_ (.I(\t2pre[8] ),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _3155_ (.A1(_0795_),
    .A2(_0796_),
    .B1(_0798_),
    .B2(_0799_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3156_ (.A1(_0778_),
    .A2(_0797_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3157_ (.A1(\t2pre[8] ),
    .A2(_0801_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3158_ (.A1(_0792_),
    .A2(_0794_),
    .A3(_0800_),
    .A4(_0802_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3159_ (.A1(_0763_),
    .A2(_0775_),
    .A3(_0790_),
    .A4(_0803_),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3160_ (.I(_0780_),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3161_ (.A1(_0805_),
    .A2(_0781_),
    .B(_0779_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3162_ (.A1(\t2pre[7] ),
    .A2(_0797_),
    .A3(_0806_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3163_ (.A1(_0797_),
    .A2(_0806_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3164_ (.I(\t2pre[5] ),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3165_ (.I(\t2pre_counter[5] ),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3166_ (.I(\t2pre_counter[4] ),
    .Z(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3167_ (.A1(_0811_),
    .A2(_0780_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _3168_ (.A1(_0810_),
    .A2(_0812_),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3169_ (.A1(_0810_),
    .A2(_0811_),
    .A3(_0805_),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3170_ (.I(\t2pre_counter[6] ),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3171_ (.A1(_0805_),
    .A2(_0781_),
    .B1(_0814_),
    .B2(_0815_),
    .C(\t2pre[6] ),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3172_ (.A1(_0809_),
    .A2(_0813_),
    .B(_0816_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3173_ (.I(\t2pre_counter[1] ),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3174_ (.I(\t2pre_counter[0] ),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3175_ (.A1(\t2pre_counter[3] ),
    .A2(\t2pre_counter[2] ),
    .A3(_0818_),
    .A4(_0819_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _3176_ (.A1(_0811_),
    .A2(_0820_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3177_ (.A1(\t2pre[4] ),
    .A2(_0821_),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3178_ (.A1(_0809_),
    .A2(_0813_),
    .B(_0822_),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3179_ (.A1(_0810_),
    .A2(_0811_),
    .A3(_0780_),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3180_ (.A1(_0805_),
    .A2(_0781_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3181_ (.A1(\t2pre_counter[6] ),
    .A2(_0824_),
    .B(_0825_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3182_ (.A1(_2040_),
    .A2(_0808_),
    .B1(_0817_),
    .B2(_0823_),
    .C1(_0826_),
    .C2(_2023_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3183_ (.I(_0819_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3184_ (.A1(_0818_),
    .A2(_0828_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _3185_ (.A1(\t2pre_counter[2] ),
    .A2(_0829_),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3186_ (.A1(\t2pre_counter[2] ),
    .A2(_0818_),
    .A3(_0819_),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3187_ (.A1(\t2pre_counter[3] ),
    .A2(_0831_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3188_ (.A1(\t2pre[2] ),
    .A2(_0830_),
    .B1(_0832_),
    .B2(\t2pre[3] ),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3189_ (.A1(_0818_),
    .A2(_0819_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3190_ (.A1(\t2pre[1] ),
    .A2(_0834_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3191_ (.A1(\t2pre[0] ),
    .A2(_0828_),
    .B1(_0834_),
    .B2(\t2pre[1] ),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3192_ (.A1(_0835_),
    .A2(_0836_),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3193_ (.A1(_1942_),
    .A2(_0830_),
    .B1(_0835_),
    .B2(_0837_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3194_ (.A1(_0833_),
    .A2(_0838_),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3195_ (.A1(_2040_),
    .A2(_0808_),
    .B1(_0826_),
    .B2(_2023_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3196_ (.A1(_0810_),
    .A2(_0812_),
    .Z(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3197_ (.A1(\t2pre[5] ),
    .A2(_0841_),
    .B1(_0821_),
    .B2(_1984_),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3198_ (.A1(_1984_),
    .A2(_0821_),
    .B1(_0832_),
    .B2(\t2pre[3] ),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3199_ (.A1(_0807_),
    .A2(_0843_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3200_ (.A1(_0840_),
    .A2(_0817_),
    .A3(_0842_),
    .A4(_0844_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3201_ (.A1(_0807_),
    .A2(_0827_),
    .B1(_0839_),
    .B2(_0845_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _3202_ (.A1(_1947_),
    .A2(_0786_),
    .B1(_0793_),
    .B2(_1923_),
    .C(_0800_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3203_ (.A1(_0790_),
    .A2(_0847_),
    .B(_0792_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3204_ (.A1(_0763_),
    .A2(_0775_),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3205_ (.I(_0768_),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3206_ (.I(\t2pre[12] ),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3207_ (.A1(_0851_),
    .A2(_0773_),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3208_ (.A1(_0772_),
    .A2(_0852_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3209_ (.A1(_0766_),
    .A2(_0853_),
    .B(_0763_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _3210_ (.A1(_0804_),
    .A2(_0846_),
    .B1(_0848_),
    .B2(_0849_),
    .C1(_0850_),
    .C2(_0854_),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3211_ (.A1(_0763_),
    .A2(_0775_),
    .A3(_0790_),
    .A4(_0803_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3212_ (.A1(_1942_),
    .A2(_0830_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3213_ (.A1(\t2pre[0] ),
    .A2(_0828_),
    .B(_0857_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3214_ (.A1(_0833_),
    .A2(_0837_),
    .A3(_0858_),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3215_ (.A1(_0787_),
    .A2(_0776_),
    .A3(_0777_),
    .A4(_0782_),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3216_ (.A1(\t2pre_counter[15] ),
    .A2(\t2pre_counter[14] ),
    .A3(_0744_),
    .A4(_0860_),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _3217_ (.A1(_0856_),
    .A2(_0845_),
    .A3(_0859_),
    .B(_0861_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3218_ (.I(\t2_top[15] ),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3219_ (.I(\timer2[15] ),
    .Z(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3220_ (.I(\timer2[14] ),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3221_ (.I(\timer2[13] ),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3222_ (.A1(\t2_top[14] ),
    .A2(_0865_),
    .B1(_0866_),
    .B2(\t2_top[13] ),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3223_ (.I(_0867_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3224_ (.I(\timer2[12] ),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3225_ (.I(\timer2[11] ),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3226_ (.A1(\t2_top[12] ),
    .A2(_0869_),
    .B1(_0870_),
    .B2(\t2_top[11] ),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3227_ (.I(\t2_top[9] ),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3228_ (.I(\timer2[9] ),
    .Z(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3229_ (.I(\timer2[8] ),
    .Z(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3230_ (.I(\t2_top[8] ),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3231_ (.A1(_0872_),
    .A2(_0873_),
    .B1(_0874_),
    .B2(_0875_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3232_ (.I(\t2_top[10] ),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _3233_ (.A1(_0877_),
    .A2(\timer2[10] ),
    .B1(\timer2[9] ),
    .B2(_0872_),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3234_ (.I(\t2_top[11] ),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3235_ (.A1(_0879_),
    .A2(\timer2[11] ),
    .B1(\timer2[10] ),
    .B2(_0877_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3236_ (.A1(_0876_),
    .A2(_0878_),
    .B(_0880_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3237_ (.I(_0866_),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3238_ (.I(_0869_),
    .Z(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3239_ (.A1(_2016_),
    .A2(_0882_),
    .B1(_0883_),
    .B2(_1998_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3240_ (.A1(_0871_),
    .A2(_0881_),
    .B(_0884_),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3241_ (.I(\timer2[14] ),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3242_ (.I(\t2_top[14] ),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3243_ (.A1(_0863_),
    .A2(_0864_),
    .B1(_0886_),
    .B2(_0887_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3244_ (.A1(_0868_),
    .A2(_0885_),
    .B(_0888_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3245_ (.A1(_0863_),
    .A2(_0864_),
    .B(_0889_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3246_ (.I(\t2_top[7] ),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3247_ (.I(\timer2[7] ),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3248_ (.I(\timer2[6] ),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3249_ (.I(\t2_top[6] ),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3250_ (.A1(_0891_),
    .A2(_0892_),
    .B1(_0893_),
    .B2(_0894_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3251_ (.I(_0895_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3252_ (.I(\t2_top[5] ),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3253_ (.I(\timer2[5] ),
    .Z(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3254_ (.I(\t2_top[4] ),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3255_ (.A1(_0897_),
    .A2(_0898_),
    .B1(\timer2[4] ),
    .B2(_0899_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3256_ (.I(\t2_top[3] ),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3257_ (.I(\timer2[3] ),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3258_ (.I(\t2_top[2] ),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3259_ (.A1(_0901_),
    .A2(_0902_),
    .B1(\timer2[2] ),
    .B2(_0903_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3260_ (.I(_0904_),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3261_ (.I(\timer2[2] ),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3262_ (.I(\t2_top[1] ),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3263_ (.I(\timer2[1] ),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3264_ (.A1(_0907_),
    .A2(_0908_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3265_ (.I(\t2_top[0] ),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3266_ (.I(\timer2[0] ),
    .Z(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3267_ (.A1(\t2_top[1] ),
    .A2(\timer2[1] ),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3268_ (.A1(_0910_),
    .A2(_0911_),
    .B(_0912_),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3269_ (.A1(\t2_top[2] ),
    .A2(_0906_),
    .B1(_0909_),
    .B2(_0913_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3270_ (.I(\timer2[4] ),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3271_ (.I(_0902_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3272_ (.A1(\t2_top[4] ),
    .A2(_0915_),
    .B1(_0916_),
    .B2(\t2_top[3] ),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3273_ (.A1(_0905_),
    .A2(_0914_),
    .B(_0917_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3274_ (.I(\timer2[5] ),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3275_ (.A1(\t2_top[5] ),
    .A2(_0919_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3276_ (.I(\timer2[6] ),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3277_ (.A1(\t2_top[6] ),
    .A2(_0921_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3278_ (.A1(_0920_),
    .A2(_0922_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3279_ (.A1(_0900_),
    .A2(_0918_),
    .B(_0923_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3280_ (.I(\timer2[7] ),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3281_ (.A1(\t2_top[7] ),
    .A2(_0925_),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3282_ (.I(_0888_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _3283_ (.A1(_2016_),
    .A2(_0882_),
    .B1(_0883_),
    .B2(_1998_),
    .C(_0880_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3284_ (.I(\timer2[15] ),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3285_ (.I(\timer2[8] ),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3286_ (.A1(\t2_top[15] ),
    .A2(_0929_),
    .B1(_0930_),
    .B2(\t2_top[8] ),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3287_ (.A1(_0867_),
    .A2(_0871_),
    .A3(_0876_),
    .A4(_0931_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3288_ (.A1(_0927_),
    .A2(_0878_),
    .A3(_0928_),
    .A4(_0932_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3289_ (.A1(_0896_),
    .A2(_0924_),
    .B(_0926_),
    .C(_0933_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3290_ (.I(\timer2[2] ),
    .Z(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3291_ (.A1(_0903_),
    .A2(_0935_),
    .B(_0920_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3292_ (.A1(_0900_),
    .A2(_0917_),
    .A3(_0904_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3293_ (.A1(_0910_),
    .A2(_0911_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3294_ (.A1(_0895_),
    .A2(_0922_),
    .A3(_0926_),
    .A4(_0938_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3295_ (.A1(_0913_),
    .A2(_0936_),
    .A3(_0937_),
    .A4(_0939_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3296_ (.A1(_0890_),
    .A2(_0934_),
    .B1(_0940_),
    .B2(_0933_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3297_ (.A1(_0855_),
    .A2(_0862_),
    .B(_0941_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3298_ (.I(_0942_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3299_ (.I(_0717_),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _3300_ (.A1(_0944_),
    .A2(_0720_),
    .B1(_0943_),
    .B2(\settings[2] ),
    .C(_0465_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3301_ (.A1(_0741_),
    .A2(_0943_),
    .B(_0945_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3302_ (.I(_0467_),
    .Z(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3303_ (.A1(_0946_),
    .A2(net18),
    .Z(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3304_ (.I(_0947_),
    .Z(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3305_ (.A1(_0946_),
    .A2(net19),
    .Z(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3306_ (.I(_0948_),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3307_ (.I(_1830_),
    .Z(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3308_ (.I(_0458_),
    .Z(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3309_ (.A1(_0949_),
    .A2(_1846_),
    .A3(_0950_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3310_ (.I(_0951_),
    .Z(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3311_ (.I(_0952_),
    .Z(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3312_ (.I(_0396_),
    .Z(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3313_ (.I(_0454_),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3314_ (.I(_0951_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3315_ (.A1(_0954_),
    .A2(_0955_),
    .B(_0956_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3316_ (.I(\timer0[0] ),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3317_ (.I(_0395_),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3318_ (.A1(_0958_),
    .A2(_0959_),
    .Z(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3319_ (.A1(\temp[0] ),
    .A2(_0953_),
    .B1(_0957_),
    .B2(_0960_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3320_ (.A1(_1785_),
    .A2(_0961_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3321_ (.I(\temp[1] ),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3322_ (.I(_0952_),
    .Z(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3323_ (.A1(_0962_),
    .A2(_0963_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3324_ (.I(_0951_),
    .Z(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3325_ (.A1(\timer0[1] ),
    .A2(_0958_),
    .A3(_0959_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3326_ (.I(_0395_),
    .Z(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3327_ (.A1(_0958_),
    .A2(_0967_),
    .B(\timer0[1] ),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _3328_ (.A1(_0455_),
    .A2(_0965_),
    .A3(_0966_),
    .A4(_0968_),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3329_ (.I(_1784_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3330_ (.A1(_0964_),
    .A2(_0969_),
    .B(_0970_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3331_ (.A1(\timer0[2] ),
    .A2(\timer0[1] ),
    .A3(_0958_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3332_ (.A1(_0955_),
    .A2(_0971_),
    .B(_0967_),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3333_ (.I(_0719_),
    .Z(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3334_ (.A1(_1898_),
    .A2(_0973_),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3335_ (.A1(\timer0[2] ),
    .A2(_0966_),
    .B(_0972_),
    .C(_0974_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3336_ (.I(\temp[2] ),
    .Z(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3337_ (.I(_0952_),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3338_ (.A1(_0976_),
    .A2(_0977_),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3339_ (.A1(_0975_),
    .A2(_0978_),
    .B(_0970_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3340_ (.I(\temp[3] ),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3341_ (.I(_0979_),
    .Z(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3342_ (.I(_0965_),
    .Z(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3343_ (.A1(_0385_),
    .A2(_0391_),
    .B(_0394_),
    .C(_0454_),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3344_ (.I(_0982_),
    .Z(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3345_ (.A1(_0406_),
    .A2(_0971_),
    .A3(_0983_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3346_ (.I(_0952_),
    .Z(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3347_ (.A1(\timer0[3] ),
    .A2(_0972_),
    .B(_0985_),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3348_ (.I(_1779_),
    .Z(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3349_ (.I(_0987_),
    .Z(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3350_ (.A1(_0980_),
    .A2(_0981_),
    .B1(_0984_),
    .B2(_0986_),
    .C(_0988_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3351_ (.I(\temp[4] ),
    .Z(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3352_ (.A1(_0989_),
    .A2(_0963_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3353_ (.I(_0395_),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3354_ (.A1(\timer0[3] ),
    .A2(_0991_),
    .A3(_0971_),
    .Z(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3355_ (.I(_0454_),
    .Z(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3356_ (.A1(\timer0[4] ),
    .A2(\timer0[3] ),
    .A3(_0971_),
    .Z(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3357_ (.A1(_0993_),
    .A2(_0994_),
    .B(_0967_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3358_ (.A1(\timer0[4] ),
    .A2(_0992_),
    .B(_0995_),
    .C(_0974_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3359_ (.A1(_0990_),
    .A2(_0996_),
    .B(_0970_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3360_ (.I(\temp[5] ),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3361_ (.A1(_0402_),
    .A2(_0983_),
    .A3(_0994_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3362_ (.A1(\timer0[5] ),
    .A2(_0995_),
    .B(_0985_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3363_ (.A1(_0997_),
    .A2(_0981_),
    .B1(_0998_),
    .B2(_0999_),
    .C(_0988_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3364_ (.I(\temp[6] ),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3365_ (.I(_1000_),
    .Z(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3366_ (.A1(\timer0[5] ),
    .A2(_0994_),
    .Z(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3367_ (.A1(_0401_),
    .A2(_0983_),
    .A3(_1002_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3368_ (.A1(_0955_),
    .A2(_1002_),
    .B(_0954_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3369_ (.A1(_0399_),
    .A2(_1004_),
    .B(_0985_),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3370_ (.I(_1779_),
    .Z(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3371_ (.I(_1006_),
    .Z(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3372_ (.A1(_1001_),
    .A2(_0977_),
    .B1(_1003_),
    .B2(_1005_),
    .C(_1007_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3373_ (.I(\temp[7] ),
    .Z(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3374_ (.A1(_1008_),
    .A2(_0953_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3375_ (.A1(_0399_),
    .A2(_1002_),
    .Z(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3376_ (.A1(_0398_),
    .A2(_0396_),
    .A3(_1010_),
    .Z(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3377_ (.A1(_0991_),
    .A2(_1010_),
    .B(_0398_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _3378_ (.A1(_0455_),
    .A2(_0965_),
    .A3(_1011_),
    .A4(_1012_),
    .Z(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3379_ (.A1(_1009_),
    .A2(_1013_),
    .B(_0970_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3380_ (.A1(\timer0[8] ),
    .A2(\timer0[7] ),
    .A3(_0399_),
    .A4(_1002_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3381_ (.A1(_0993_),
    .A2(_1014_),
    .B(_0967_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3382_ (.A1(\timer0[8] ),
    .A2(_1011_),
    .B(_1015_),
    .C(_0974_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3383_ (.A1(_0724_),
    .A2(_0963_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3384_ (.I(_1780_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3385_ (.I(_1018_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3386_ (.A1(_1016_),
    .A2(_1017_),
    .B(_1019_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3387_ (.I(_0728_),
    .Z(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3388_ (.A1(_0423_),
    .A2(_0983_),
    .A3(_1014_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3389_ (.A1(\timer0[9] ),
    .A2(_1015_),
    .B(_0985_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3390_ (.A1(_1020_),
    .A2(_0977_),
    .B1(_1021_),
    .B2(_1022_),
    .C(_1007_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3391_ (.I(_0731_),
    .Z(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3392_ (.A1(\timer0[9] ),
    .A2(_1014_),
    .Z(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3393_ (.A1(_0427_),
    .A2(_0982_),
    .A3(_1024_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3394_ (.A1(_0955_),
    .A2(_1024_),
    .B(_0991_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3395_ (.A1(_0420_),
    .A2(_1026_),
    .B(_0965_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3396_ (.A1(_1023_),
    .A2(_0977_),
    .B1(_1025_),
    .B2(_1027_),
    .C(_1007_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3397_ (.I(_0457_),
    .Z(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3398_ (.A1(_1028_),
    .A2(_0953_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3399_ (.I(\timer0[11] ),
    .Z(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3400_ (.A1(_0420_),
    .A2(_1024_),
    .Z(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3401_ (.A1(_1030_),
    .A2(_0396_),
    .A3(_1031_),
    .Z(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3402_ (.A1(_0991_),
    .A2(_1031_),
    .B(_1030_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _3403_ (.A1(_0455_),
    .A2(_0956_),
    .A3(_1032_),
    .A4(_1033_),
    .Z(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3404_ (.A1(_1029_),
    .A2(_1034_),
    .B(_1019_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3405_ (.A1(\timer0[12] ),
    .A2(_1030_),
    .A3(_0420_),
    .A4(_1024_),
    .Z(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3406_ (.A1(_0993_),
    .A2(_1035_),
    .B(_0959_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3407_ (.A1(\timer0[12] ),
    .A2(_1032_),
    .B(_1036_),
    .C(_0974_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3408_ (.I(net13),
    .Z(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3409_ (.I(_1038_),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3410_ (.A1(_1039_),
    .A2(_0963_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3411_ (.A1(_1037_),
    .A2(_1040_),
    .B(_1019_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3412_ (.I(_0944_),
    .Z(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3413_ (.A1(_0436_),
    .A2(_1035_),
    .Z(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3414_ (.A1(\timer0[13] ),
    .A2(_1036_),
    .B1(_1042_),
    .B2(_0982_),
    .C(_0956_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3415_ (.I(_1783_),
    .Z(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3416_ (.I(_1044_),
    .Z(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3417_ (.A1(_1041_),
    .A2(_0981_),
    .B(_1043_),
    .C(_1045_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3418_ (.I(_0735_),
    .Z(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3419_ (.A1(\timer0[13] ),
    .A2(_1035_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3420_ (.A1(_0439_),
    .A2(_1047_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3421_ (.I(_1047_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3422_ (.A1(_0993_),
    .A2(_1049_),
    .B(_0959_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3423_ (.A1(_0982_),
    .A2(_1048_),
    .B1(_1050_),
    .B2(_0439_),
    .C(_0956_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3424_ (.A1(_1046_),
    .A2(_0981_),
    .B(_1051_),
    .C(_1045_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3425_ (.I(net16),
    .Z(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3426_ (.A1(_1052_),
    .A2(_0953_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3427_ (.A1(_0439_),
    .A2(_0954_),
    .A3(_1049_),
    .Z(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3428_ (.A1(\timer0[15] ),
    .A2(_1054_),
    .B(_0957_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3429_ (.A1(_1053_),
    .A2(_1055_),
    .B(_1019_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3430_ (.I(\temp[0] ),
    .Z(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3431_ (.A1(_1841_),
    .A2(_1854_),
    .A3(_0950_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3432_ (.I(_1057_),
    .Z(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3433_ (.I(_1058_),
    .Z(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3434_ (.A1(_1056_),
    .A2(_1059_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3435_ (.I(_0642_),
    .Z(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3436_ (.I(_0718_),
    .Z(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3437_ (.A1(_1843_),
    .A2(_1062_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3438_ (.I(_1063_),
    .Z(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3439_ (.I(\timer1[0] ),
    .Z(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3440_ (.A1(_0574_),
    .A2(_0583_),
    .B(_0473_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3441_ (.A1(_1065_),
    .A2(_1066_),
    .Z(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3442_ (.A1(_1061_),
    .A2(_1064_),
    .A3(_1067_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3443_ (.I(_1018_),
    .Z(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3444_ (.A1(_1060_),
    .A2(_1068_),
    .B(_1069_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3445_ (.A1(_0962_),
    .A2(_1059_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3446_ (.I(_1066_),
    .Z(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3447_ (.A1(_0617_),
    .A2(_1065_),
    .A3(_1071_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3448_ (.I(\timer1[0] ),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3449_ (.I(_0473_),
    .Z(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3450_ (.I(_1074_),
    .Z(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3451_ (.I(_0584_),
    .Z(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3452_ (.I(_1076_),
    .Z(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3453_ (.A1(_1073_),
    .A2(_1075_),
    .A3(_1077_),
    .B(_0615_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3454_ (.A1(_1061_),
    .A2(_1064_),
    .A3(_1072_),
    .A4(_1078_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3455_ (.A1(_1070_),
    .A2(_1079_),
    .B(_1069_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3456_ (.I(_1066_),
    .Z(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3457_ (.A1(_0617_),
    .A2(_1065_),
    .A3(_1080_),
    .Z(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3458_ (.I(_0641_),
    .Z(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3459_ (.I(_1082_),
    .Z(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3460_ (.A1(\timer1[2] ),
    .A2(_0617_),
    .A3(_1065_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3461_ (.A1(_1083_),
    .A2(_1084_),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3462_ (.A1(_1074_),
    .A2(_1076_),
    .Z(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3463_ (.I(_1086_),
    .Z(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3464_ (.I(_1063_),
    .Z(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _3465_ (.A1(\timer1[2] ),
    .A2(_1081_),
    .B1(_1085_),
    .B2(_1087_),
    .C(_1088_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3466_ (.I(_1058_),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3467_ (.A1(_0976_),
    .A2(_1090_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3468_ (.A1(_1089_),
    .A2(_1091_),
    .B(_1069_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3469_ (.I(_1057_),
    .Z(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3470_ (.I(_1092_),
    .Z(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3471_ (.I(\timer1[3] ),
    .Z(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3472_ (.A1(_1087_),
    .A2(_1085_),
    .B(_1094_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3473_ (.A1(_1066_),
    .A2(_0641_),
    .Z(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3474_ (.I(_1096_),
    .Z(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3475_ (.A1(_1094_),
    .A2(_1084_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3476_ (.I(_1058_),
    .Z(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3477_ (.A1(_1097_),
    .A2(_1098_),
    .B(_1099_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3478_ (.A1(_0980_),
    .A2(_1093_),
    .B1(_1095_),
    .B2(_1100_),
    .C(_1007_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3479_ (.I(_1058_),
    .Z(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3480_ (.A1(\temp[4] ),
    .A2(_1101_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3481_ (.A1(_0614_),
    .A2(_0615_),
    .A3(_1073_),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3482_ (.A1(_1094_),
    .A2(_1080_),
    .A3(_1103_),
    .Z(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3483_ (.A1(_0626_),
    .A2(_1094_),
    .A3(_1103_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3484_ (.A1(_1083_),
    .A2(_1105_),
    .Z(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _3485_ (.A1(_0626_),
    .A2(_1104_),
    .B1(_1106_),
    .B2(_1087_),
    .C(_1088_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3486_ (.A1(_1102_),
    .A2(_1107_),
    .B(_1069_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3487_ (.I(_1086_),
    .Z(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3488_ (.A1(_1108_),
    .A2(_1106_),
    .B(\timer1[5] ),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3489_ (.A1(\timer1[5] ),
    .A2(_1105_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3490_ (.A1(_1097_),
    .A2(_1110_),
    .B(_1099_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3491_ (.I(_1006_),
    .Z(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3492_ (.A1(_0997_),
    .A2(_1093_),
    .B1(_1109_),
    .B2(_1111_),
    .C(_1112_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3493_ (.A1(_0628_),
    .A2(_1105_),
    .Z(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3494_ (.A1(_1083_),
    .A2(_1113_),
    .Z(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3495_ (.I(\timer1[6] ),
    .Z(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3496_ (.A1(_1108_),
    .A2(_1114_),
    .B(_1115_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3497_ (.A1(_1115_),
    .A2(_1113_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3498_ (.A1(_1097_),
    .A2(_1117_),
    .B(_1099_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3499_ (.A1(_1001_),
    .A2(_1093_),
    .B1(_1116_),
    .B2(_1118_),
    .C(_1112_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3500_ (.A1(_1008_),
    .A2(_1101_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3501_ (.A1(_0628_),
    .A2(_1105_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3502_ (.A1(\timer1[7] ),
    .A2(_1115_),
    .A3(_1071_),
    .A4(_1120_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3503_ (.I(_1076_),
    .Z(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3504_ (.A1(_1115_),
    .A2(_1120_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3505_ (.A1(_1075_),
    .A2(_1122_),
    .A3(_1123_),
    .B(_0631_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3506_ (.A1(_1061_),
    .A2(_1064_),
    .A3(_1121_),
    .A4(_1124_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3507_ (.I(_1018_),
    .Z(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3508_ (.A1(_1119_),
    .A2(_1125_),
    .B(_1126_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3509_ (.I(_1074_),
    .Z(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3510_ (.I(_1076_),
    .Z(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _3511_ (.A1(_0631_),
    .A2(_1127_),
    .A3(_1128_),
    .A4(_1123_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3512_ (.A1(\timer1[8] ),
    .A2(\timer1[7] ),
    .A3(\timer1[6] ),
    .A4(_1120_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3513_ (.A1(_1082_),
    .A2(_1130_),
    .Z(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _3514_ (.A1(\timer1[8] ),
    .A2(_1129_),
    .B1(_1131_),
    .B2(_1087_),
    .C(_1063_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3515_ (.A1(_0724_),
    .A2(_1059_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3516_ (.A1(_1132_),
    .A2(_1133_),
    .B(_1126_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3517_ (.A1(_1108_),
    .A2(_1131_),
    .B(\timer1[9] ),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3518_ (.A1(\timer1[9] ),
    .A2(_1130_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3519_ (.A1(_1097_),
    .A2(_1135_),
    .B(_1092_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3520_ (.A1(_1020_),
    .A2(_1090_),
    .B1(_1134_),
    .B2(_1136_),
    .C(_1112_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3521_ (.A1(_0596_),
    .A2(_1130_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3522_ (.A1(_0600_),
    .A2(_1096_),
    .A3(_1137_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3523_ (.A1(_0596_),
    .A2(_1130_),
    .B(_1082_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3524_ (.A1(_1080_),
    .A2(_1139_),
    .B(_0600_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3525_ (.A1(_1099_),
    .A2(_1140_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3526_ (.A1(_1023_),
    .A2(_1090_),
    .B1(_1138_),
    .B2(_1141_),
    .C(_1112_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3527_ (.I(net12),
    .Z(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3528_ (.A1(_1142_),
    .A2(_1101_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3529_ (.A1(\timer1[11] ),
    .A2(\timer1[10] ),
    .A3(_1071_),
    .A4(_1137_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3530_ (.A1(\timer1[10] ),
    .A2(_1137_),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3531_ (.A1(_1127_),
    .A2(_1122_),
    .A3(_1145_),
    .B(_0602_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3532_ (.A1(_1061_),
    .A2(_1064_),
    .A3(_1144_),
    .A4(_1146_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3533_ (.A1(_1143_),
    .A2(_1147_),
    .B(_1126_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _3534_ (.A1(_0602_),
    .A2(_1127_),
    .A3(_1122_),
    .A4(_1145_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3535_ (.A1(_0592_),
    .A2(\timer1[11] ),
    .A3(\timer1[10] ),
    .A4(_1137_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3536_ (.A1(_1082_),
    .A2(_1149_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3537_ (.A1(_1080_),
    .A2(_1150_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3538_ (.A1(_0592_),
    .A2(_1148_),
    .B(_1151_),
    .C(_1088_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3539_ (.A1(_1039_),
    .A2(_1059_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3540_ (.A1(_1152_),
    .A2(_1153_),
    .B(_1126_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3541_ (.A1(\timer1[13] ),
    .A2(_1149_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3542_ (.A1(\timer1[13] ),
    .A2(_1151_),
    .B1(_1154_),
    .B2(_1096_),
    .C(_1092_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3543_ (.A1(_1041_),
    .A2(_1093_),
    .B(_1155_),
    .C(_1045_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3544_ (.A1(_0589_),
    .A2(_1149_),
    .Z(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3545_ (.A1(_1083_),
    .A2(_1156_),
    .Z(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3546_ (.A1(_1108_),
    .A2(_1157_),
    .B(_0588_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3547_ (.A1(_0588_),
    .A2(_1156_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3548_ (.A1(_1096_),
    .A2(_1159_),
    .B(_1092_),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3549_ (.I(_1006_),
    .Z(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3550_ (.A1(_0735_),
    .A2(_1090_),
    .B1(_1158_),
    .B2(_1160_),
    .C(_1161_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3551_ (.A1(_1052_),
    .A2(_1101_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _3552_ (.A1(_0635_),
    .A2(_1127_),
    .A3(_1122_),
    .A4(_1156_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3553_ (.A1(\timer1[15] ),
    .A2(_1163_),
    .B(_1088_),
    .C(_0642_),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3554_ (.I(_1018_),
    .Z(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3555_ (.A1(_1162_),
    .A2(_1164_),
    .B(_1165_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3556_ (.A1(_1859_),
    .A2(_1822_),
    .A3(_0459_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3557_ (.I(_1166_),
    .Z(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3558_ (.I(_1167_),
    .Z(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3559_ (.I(_1168_),
    .Z(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3560_ (.I(_1166_),
    .Z(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3561_ (.I(_1170_),
    .Z(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3562_ (.A1(\t0_capture[0] ),
    .A2(_1171_),
    .B(_0733_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3563_ (.A1(_0409_),
    .A2(_1169_),
    .B(_1172_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3564_ (.A1(\t0_capture[1] ),
    .A2(_1171_),
    .B(_0733_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3565_ (.A1(_0408_),
    .A2(_1169_),
    .B(_1173_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3566_ (.I(_1804_),
    .Z(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3567_ (.A1(\t0_capture[2] ),
    .A2(_1171_),
    .B(_1174_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3568_ (.A1(_0411_),
    .A2(_1169_),
    .B(_1175_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3569_ (.A1(\t0_capture[3] ),
    .A2(_1171_),
    .B(_1174_),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3570_ (.A1(_0406_),
    .A2(_1169_),
    .B(_1176_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3571_ (.I(_1168_),
    .Z(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3572_ (.I(_1170_),
    .Z(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3573_ (.A1(\t0_capture[4] ),
    .A2(_1178_),
    .B(_1174_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3574_ (.A1(_0405_),
    .A2(_1177_),
    .B(_1179_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3575_ (.A1(\t0_capture[5] ),
    .A2(_1178_),
    .B(_1174_),
    .ZN(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3576_ (.A1(_0402_),
    .A2(_1177_),
    .B(_1180_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3577_ (.I(_1803_),
    .Z(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3578_ (.I(_1181_),
    .Z(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3579_ (.A1(\t0_capture[6] ),
    .A2(_1178_),
    .B(_1182_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3580_ (.A1(_0401_),
    .A2(_1177_),
    .B(_1183_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3581_ (.I(_0398_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3582_ (.A1(\t0_capture[7] ),
    .A2(_1178_),
    .B(_1182_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3583_ (.A1(_1184_),
    .A2(_1177_),
    .B(_1185_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3584_ (.I(_1167_),
    .Z(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3585_ (.I(_1186_),
    .Z(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3586_ (.I(_1167_),
    .Z(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3587_ (.I(_1188_),
    .Z(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3588_ (.A1(\t0_capture[8] ),
    .A2(_1189_),
    .B(_1182_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3589_ (.A1(_0424_),
    .A2(_1187_),
    .B(_1190_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3590_ (.A1(\t0_capture[9] ),
    .A2(_1189_),
    .B(_1182_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3591_ (.A1(_0423_),
    .A2(_1187_),
    .B(_1191_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3592_ (.I(_1181_),
    .Z(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3593_ (.A1(\t0_capture[10] ),
    .A2(_1189_),
    .B(_1192_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3594_ (.A1(_0427_),
    .A2(_1187_),
    .B(_1193_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3595_ (.A1(_1864_),
    .A2(_1815_),
    .A3(_1062_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3596_ (.I(_1194_),
    .Z(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3597_ (.A1(\t0_capture[11] ),
    .A2(_1195_),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3598_ (.I(_1170_),
    .Z(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3599_ (.A1(_1030_),
    .A2(_1197_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3600_ (.A1(_1196_),
    .A2(_1198_),
    .B(_1165_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3601_ (.A1(\t0_capture[12] ),
    .A2(_1189_),
    .B(_1192_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3602_ (.A1(_0442_),
    .A2(_1187_),
    .B(_1199_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3603_ (.I(_1186_),
    .Z(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3604_ (.I(_1188_),
    .Z(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3605_ (.A1(\t0_capture[13] ),
    .A2(_1201_),
    .B(_1192_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3606_ (.A1(_0436_),
    .A2(_1200_),
    .B(_1202_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3607_ (.A1(\t0_capture[14] ),
    .A2(_1201_),
    .B(_1192_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3608_ (.A1(_0431_),
    .A2(_1200_),
    .B(_1203_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3609_ (.I(_1181_),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3610_ (.A1(\t0_capture[15] ),
    .A2(_1201_),
    .B(_1204_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3611_ (.A1(_0434_),
    .A2(_1200_),
    .B(_1205_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3612_ (.A1(\t1_capture[0] ),
    .A2(_1201_),
    .B(_1204_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3613_ (.A1(_1073_),
    .A2(_1200_),
    .B(_1206_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3614_ (.I(_1186_),
    .Z(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3615_ (.I(_1188_),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3616_ (.A1(\t1_capture[1] ),
    .A2(_1208_),
    .B(_1204_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3617_ (.A1(_0615_),
    .A2(_1207_),
    .B(_1209_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3618_ (.A1(\t1_capture[2] ),
    .A2(_1208_),
    .B(_1204_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3619_ (.A1(_0614_),
    .A2(_1207_),
    .B(_1210_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3620_ (.I(_1181_),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3621_ (.A1(\t1_capture[3] ),
    .A2(_1208_),
    .B(_1211_),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3622_ (.A1(_0621_),
    .A2(_1207_),
    .B(_1212_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3623_ (.A1(\t1_capture[4] ),
    .A2(_1195_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3624_ (.A1(_0626_),
    .A2(_1197_),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3625_ (.A1(_1213_),
    .A2(_1214_),
    .B(_1165_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3626_ (.A1(\t1_capture[5] ),
    .A2(_1208_),
    .B(_1211_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3627_ (.A1(_0628_),
    .A2(_1207_),
    .B(_1215_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3628_ (.I(_1186_),
    .Z(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3629_ (.I(_1188_),
    .Z(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3630_ (.A1(\t1_capture[6] ),
    .A2(_1217_),
    .B(_1211_),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3631_ (.A1(_0612_),
    .A2(_1216_),
    .B(_1218_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3632_ (.A1(\t1_capture[7] ),
    .A2(_1217_),
    .B(_1211_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3633_ (.A1(_0631_),
    .A2(_1216_),
    .B(_1219_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3634_ (.I(_1803_),
    .Z(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3635_ (.I(_1220_),
    .Z(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3636_ (.A1(\t1_capture[8] ),
    .A2(_1217_),
    .B(_1221_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3637_ (.A1(_0597_),
    .A2(_1216_),
    .B(_1222_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3638_ (.A1(\t1_capture[9] ),
    .A2(_1217_),
    .B(_1221_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3639_ (.A1(_0596_),
    .A2(_1216_),
    .B(_1223_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3640_ (.I(_1167_),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3641_ (.I(_1224_),
    .Z(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3642_ (.I(_1166_),
    .Z(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3643_ (.I(_1226_),
    .Z(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3644_ (.A1(\t1_capture[10] ),
    .A2(_1227_),
    .B(_1221_),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3645_ (.A1(_0600_),
    .A2(_1225_),
    .B(_1228_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3646_ (.A1(\t1_capture[11] ),
    .A2(_1227_),
    .B(_1221_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3647_ (.A1(_0602_),
    .A2(_1225_),
    .B(_1229_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3648_ (.A1(\t1_capture[12] ),
    .A2(_1195_),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3649_ (.I(_1170_),
    .Z(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3650_ (.A1(_0592_),
    .A2(_1231_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3651_ (.A1(_1230_),
    .A2(_1232_),
    .B(_1165_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3652_ (.I(_1220_),
    .Z(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3653_ (.A1(\t1_capture[13] ),
    .A2(_1227_),
    .B(_1233_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3654_ (.A1(_0589_),
    .A2(_1225_),
    .B(_1234_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3655_ (.A1(\t1_capture[14] ),
    .A2(_1227_),
    .B(_1233_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3656_ (.A1(_0635_),
    .A2(_1225_),
    .B(_1235_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3657_ (.I(_1224_),
    .Z(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3658_ (.I(_1226_),
    .Z(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3659_ (.A1(\t1_capture[15] ),
    .A2(_1237_),
    .B(_1233_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3660_ (.A1(_0585_),
    .A2(_1236_),
    .B(_1238_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3661_ (.I(_0911_),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3662_ (.I(_1239_),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3663_ (.A1(\t2_capture[0] ),
    .A2(_1237_),
    .B(_1233_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3664_ (.A1(_1240_),
    .A2(_1236_),
    .B(_1241_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3665_ (.A1(\t2_capture[1] ),
    .A2(_1195_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3666_ (.I(_0908_),
    .Z(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3667_ (.A1(_1243_),
    .A2(_1231_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3668_ (.I(_1783_),
    .Z(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3669_ (.I(_1245_),
    .Z(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3670_ (.A1(_1242_),
    .A2(_1244_),
    .B(_1246_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3671_ (.I(_1220_),
    .Z(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3672_ (.A1(\t2_capture[2] ),
    .A2(_1237_),
    .B(_1247_),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3673_ (.A1(_0906_),
    .A2(_1236_),
    .B(_1248_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3674_ (.A1(\t2_capture[3] ),
    .A2(_1237_),
    .B(_1247_),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3675_ (.A1(_0916_),
    .A2(_1236_),
    .B(_1249_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3676_ (.I(_1224_),
    .Z(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3677_ (.I(_1226_),
    .Z(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3678_ (.A1(\t2_capture[4] ),
    .A2(_1251_),
    .B(_1247_),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3679_ (.A1(_0915_),
    .A2(_1250_),
    .B(_1252_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3680_ (.A1(\t2_capture[5] ),
    .A2(_1251_),
    .B(_1247_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3681_ (.A1(_0919_),
    .A2(_1250_),
    .B(_1253_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3682_ (.I(_1220_),
    .Z(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3683_ (.A1(\t2_capture[6] ),
    .A2(_1251_),
    .B(_1254_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3684_ (.A1(_0921_),
    .A2(_1250_),
    .B(_1255_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3685_ (.A1(\t2_capture[7] ),
    .A2(_1251_),
    .B(_1254_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3686_ (.A1(_0925_),
    .A2(_1250_),
    .B(_1256_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3687_ (.I(_1224_),
    .Z(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3688_ (.I(_1226_),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3689_ (.A1(\t2_capture[8] ),
    .A2(_1258_),
    .B(_1254_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3690_ (.A1(_0930_),
    .A2(_1257_),
    .B(_1259_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3691_ (.A1(\t2_capture[9] ),
    .A2(_1194_),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3692_ (.I(_0873_),
    .Z(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3693_ (.A1(_1261_),
    .A2(_1231_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3694_ (.A1(_1260_),
    .A2(_1262_),
    .B(_1246_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3695_ (.A1(\t2_capture[10] ),
    .A2(_1194_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3696_ (.I(\timer2[10] ),
    .Z(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3697_ (.A1(_1264_),
    .A2(_1231_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3698_ (.A1(_1263_),
    .A2(_1265_),
    .B(_1246_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3699_ (.A1(\t2_capture[11] ),
    .A2(_1258_),
    .B(_1254_),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3700_ (.A1(_0870_),
    .A2(_1257_),
    .B(_1266_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3701_ (.I(_0463_),
    .Z(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3702_ (.I(_1267_),
    .Z(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3703_ (.A1(\t2_capture[12] ),
    .A2(_1258_),
    .B(_1268_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3704_ (.A1(_0883_),
    .A2(_1257_),
    .B(_1269_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3705_ (.A1(\t2_capture[13] ),
    .A2(_1258_),
    .B(_1268_),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3706_ (.A1(_0882_),
    .A2(_1257_),
    .B(_1270_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3707_ (.A1(\t2_capture[14] ),
    .A2(_1168_),
    .B(_1268_),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3708_ (.A1(_0865_),
    .A2(_1197_),
    .B(_1271_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3709_ (.A1(\t2_capture[15] ),
    .A2(_1168_),
    .B(_1268_),
    .ZN(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3710_ (.A1(_0929_),
    .A2(_1197_),
    .B(_1272_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3711_ (.I(_0718_),
    .Z(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3712_ (.A1(_1833_),
    .A2(_1273_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3713_ (.I(_1274_),
    .Z(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3714_ (.A1(\t0pre[0] ),
    .A2(_1275_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3715_ (.I(\temp[0] ),
    .Z(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3716_ (.I(_0459_),
    .Z(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3717_ (.A1(_0949_),
    .A2(_1822_),
    .A3(_1278_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3718_ (.I(_1279_),
    .Z(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3719_ (.I(_1280_),
    .Z(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3720_ (.A1(_1277_),
    .A2(_1281_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3721_ (.A1(_1276_),
    .A2(_1282_),
    .B(_1246_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3722_ (.I(\temp[1] ),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3723_ (.I(_1283_),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3724_ (.I(_1279_),
    .Z(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3725_ (.I(_1285_),
    .Z(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3726_ (.I(_1280_),
    .Z(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3727_ (.I(_1267_),
    .Z(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3728_ (.A1(\t0pre[1] ),
    .A2(_1287_),
    .B(_1288_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3729_ (.A1(_1284_),
    .A2(_1286_),
    .B(_1289_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _3730_ (.I(\temp[2] ),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3731_ (.A1(_1945_),
    .A2(_1287_),
    .B(_1288_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3732_ (.A1(_1290_),
    .A2(_1286_),
    .B(_1291_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3733_ (.I(_0979_),
    .Z(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3734_ (.I(_1280_),
    .Z(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3735_ (.A1(\t0pre[3] ),
    .A2(_1293_),
    .B(_1288_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3736_ (.A1(_1292_),
    .A2(_1286_),
    .B(_1294_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3737_ (.A1(_1987_),
    .A2(_1275_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3738_ (.I(\temp[4] ),
    .Z(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3739_ (.A1(_1296_),
    .A2(_1281_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3740_ (.I(_1245_),
    .Z(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3741_ (.A1(_1295_),
    .A2(_1297_),
    .B(_1298_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3742_ (.I(_0997_),
    .Z(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3743_ (.A1(_2007_),
    .A2(_1293_),
    .B(_1288_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3744_ (.A1(_1299_),
    .A2(_1286_),
    .B(_1300_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3745_ (.I(_1000_),
    .Z(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3746_ (.I(_1285_),
    .Z(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3747_ (.I(_1267_),
    .Z(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3748_ (.A1(\t0pre[6] ),
    .A2(_1293_),
    .B(_1303_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3749_ (.A1(_1301_),
    .A2(_1302_),
    .B(_1304_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3750_ (.I(\temp[7] ),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3751_ (.I(_1305_),
    .Z(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3752_ (.A1(\t0pre[7] ),
    .A2(_1293_),
    .B(_1303_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3753_ (.A1(_1306_),
    .A2(_1302_),
    .B(_1307_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3754_ (.I(net9),
    .Z(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3755_ (.A1(_1308_),
    .A2(_1274_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3756_ (.A1(_0325_),
    .A2(_1275_),
    .B(_1309_),
    .C(_1045_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3757_ (.A1(\t0pre[9] ),
    .A2(_1285_),
    .B(_1303_),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3758_ (.A1(_0729_),
    .A2(_1302_),
    .B(_1310_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3759_ (.A1(\t0pre[10] ),
    .A2(_1285_),
    .B(_1303_),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3760_ (.A1(_0732_),
    .A2(_1302_),
    .B(_1311_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3761_ (.A1(_1142_),
    .A2(_1274_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3762_ (.I(_1044_),
    .Z(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3763_ (.A1(_2092_),
    .A2(_1275_),
    .B(_1312_),
    .C(_1313_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3764_ (.I(_1280_),
    .Z(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3765_ (.I(_1038_),
    .Z(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3766_ (.A1(_1315_),
    .A2(_1281_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3767_ (.I(_0463_),
    .Z(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3768_ (.I(_1317_),
    .Z(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3769_ (.I(_1318_),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3770_ (.A1(_0381_),
    .A2(_1314_),
    .B(_1316_),
    .C(_1319_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3771_ (.I(_0717_),
    .Z(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3772_ (.A1(_1320_),
    .A2(_1281_),
    .ZN(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3773_ (.A1(_2085_),
    .A2(_1314_),
    .B(_1321_),
    .C(_1319_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3774_ (.I(net15),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3775_ (.A1(_1322_),
    .A2(_1287_),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3776_ (.A1(_2058_),
    .A2(_1314_),
    .B(_1323_),
    .C(_1319_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3777_ (.I(_0738_),
    .Z(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3778_ (.A1(_1324_),
    .A2(_1287_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3779_ (.A1(_2079_),
    .A2(_1314_),
    .B(_1325_),
    .C(_1319_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3780_ (.A1(_1871_),
    .A2(_1062_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3781_ (.I(_1326_),
    .Z(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3782_ (.A1(_1895_),
    .A2(_1327_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3783_ (.A1(_1868_),
    .A2(_1869_),
    .A3(_0950_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3784_ (.I(_1329_),
    .Z(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3785_ (.I(_1330_),
    .Z(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3786_ (.A1(_1277_),
    .A2(_1331_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3787_ (.A1(_1328_),
    .A2(_1332_),
    .B(_1298_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3788_ (.I(_1330_),
    .Z(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3789_ (.I(_1329_),
    .Z(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3790_ (.I(_1267_),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3791_ (.A1(\t1pre[1] ),
    .A2(_1334_),
    .B(_1335_),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3792_ (.A1(_1284_),
    .A2(_1333_),
    .B(_1336_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3793_ (.A1(_1951_),
    .A2(_1334_),
    .B(_1335_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3794_ (.A1(_1290_),
    .A2(_1333_),
    .B(_1337_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3795_ (.A1(\t1pre[3] ),
    .A2(_1334_),
    .B(_1335_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3796_ (.A1(_1292_),
    .A2(_1333_),
    .B(_1338_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3797_ (.A1(\t1pre[4] ),
    .A2(_1327_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3798_ (.I(_1330_),
    .Z(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3799_ (.A1(_1296_),
    .A2(_1340_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3800_ (.A1(_1339_),
    .A2(_1341_),
    .B(_1298_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3801_ (.A1(_2012_),
    .A2(_1334_),
    .B(_1335_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3802_ (.A1(_1299_),
    .A2(_1333_),
    .B(_1342_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3803_ (.I(_1330_),
    .Z(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3804_ (.I(_1329_),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3805_ (.I(_0463_),
    .Z(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3806_ (.I(_1345_),
    .Z(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3807_ (.A1(_2030_),
    .A2(_1344_),
    .B(_1346_),
    .ZN(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3808_ (.A1(_1301_),
    .A2(_1343_),
    .B(_1347_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3809_ (.A1(\t1pre[7] ),
    .A2(_1344_),
    .B(_1346_),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3810_ (.A1(_1306_),
    .A2(_1343_),
    .B(_1348_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3811_ (.I(_1326_),
    .Z(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3812_ (.A1(_1308_),
    .A2(_1327_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3813_ (.A1(_0517_),
    .A2(_1349_),
    .B(_1350_),
    .C(_1313_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3814_ (.A1(_1929_),
    .A2(_1344_),
    .B(_1346_),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3815_ (.A1(_0729_),
    .A2(_1343_),
    .B(_1351_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3816_ (.A1(\t1pre[10] ),
    .A2(_1344_),
    .B(_1346_),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3817_ (.A1(_0732_),
    .A2(_1343_),
    .B(_1352_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3818_ (.A1(_1972_),
    .A2(_1327_),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3819_ (.I(_0457_),
    .Z(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3820_ (.A1(_1354_),
    .A2(_1340_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3821_ (.A1(_1353_),
    .A2(_1355_),
    .B(_1298_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3822_ (.I(_0464_),
    .Z(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3823_ (.I(_1356_),
    .Z(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3824_ (.A1(\t1pre[12] ),
    .A2(_1349_),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3825_ (.A1(_1039_),
    .A2(_1331_),
    .ZN(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3826_ (.A1(_1357_),
    .A2(_1358_),
    .A3(_1359_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3827_ (.A1(_1320_),
    .A2(_1340_),
    .ZN(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3828_ (.I(_1318_),
    .Z(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3829_ (.A1(_0491_),
    .A2(_1331_),
    .B(_1360_),
    .C(_1361_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3830_ (.A1(\t1pre[14] ),
    .A2(_1349_),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3831_ (.A1(_1046_),
    .A2(_1349_),
    .B(_1362_),
    .C(_1361_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3832_ (.A1(_1324_),
    .A2(_1340_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3833_ (.A1(_0485_),
    .A2(_1331_),
    .B(_1363_),
    .C(_1361_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3834_ (.A1(_1852_),
    .A2(_1062_),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3835_ (.I(_1364_),
    .Z(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3836_ (.A1(\t2pre[0] ),
    .A2(_1365_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3837_ (.A1(_1868_),
    .A2(_0949_),
    .A3(_0950_),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3838_ (.I(_1367_),
    .Z(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3839_ (.I(_1368_),
    .Z(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3840_ (.A1(_1277_),
    .A2(_1369_),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3841_ (.I(_1245_),
    .Z(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3842_ (.A1(_1366_),
    .A2(_1370_),
    .B(_1371_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3843_ (.I(_1368_),
    .Z(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3844_ (.I(_1367_),
    .Z(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3845_ (.I(_1345_),
    .Z(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3846_ (.A1(\t2pre[1] ),
    .A2(_1373_),
    .B(_1374_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3847_ (.A1(_1284_),
    .A2(_1372_),
    .B(_1375_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3848_ (.A1(_1942_),
    .A2(_1373_),
    .B(_1374_),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3849_ (.A1(_1290_),
    .A2(_1372_),
    .B(_1376_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3850_ (.A1(\t2pre[3] ),
    .A2(_1373_),
    .B(_1374_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3851_ (.A1(_1292_),
    .A2(_1372_),
    .B(_1377_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3852_ (.A1(_1984_),
    .A2(_1365_),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3853_ (.I(_1368_),
    .Z(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3854_ (.A1(_1296_),
    .A2(_1379_),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3855_ (.A1(_1378_),
    .A2(_1380_),
    .B(_1371_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3856_ (.A1(\t2pre[5] ),
    .A2(_1373_),
    .B(_1374_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3857_ (.A1(_1299_),
    .A2(_1372_),
    .B(_1381_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3858_ (.I(_1368_),
    .Z(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3859_ (.I(_1367_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3860_ (.I(_1345_),
    .Z(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3861_ (.A1(_2023_),
    .A2(_1383_),
    .B(_1384_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3862_ (.A1(_1301_),
    .A2(_1382_),
    .B(_1385_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3863_ (.A1(_2040_),
    .A2(_1383_),
    .B(_1384_),
    .ZN(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3864_ (.A1(_1306_),
    .A2(_1382_),
    .B(_1386_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3865_ (.I(_1364_),
    .Z(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3866_ (.A1(_0723_),
    .A2(_1365_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3867_ (.A1(_0799_),
    .A2(_1387_),
    .B(_1388_),
    .C(_1313_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3868_ (.A1(_1923_),
    .A2(_1383_),
    .B(_1384_),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3869_ (.A1(_0729_),
    .A2(_1382_),
    .B(_1389_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3870_ (.A1(_1947_),
    .A2(_1383_),
    .B(_1384_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3871_ (.A1(_0732_),
    .A2(_1382_),
    .B(_1390_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3872_ (.A1(_1142_),
    .A2(_1365_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3873_ (.A1(_0791_),
    .A2(_1387_),
    .B(_1391_),
    .C(_1313_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3874_ (.A1(_1315_),
    .A2(_1379_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3875_ (.A1(_0851_),
    .A2(_1369_),
    .B(_1392_),
    .C(_1361_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3876_ (.A1(_1320_),
    .A2(_1379_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3877_ (.I(_1318_),
    .Z(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3878_ (.A1(_0771_),
    .A2(_1369_),
    .B(_1393_),
    .C(_1394_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3879_ (.A1(\t2pre[14] ),
    .A2(_1387_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3880_ (.A1(_1046_),
    .A2(_1387_),
    .B(_1395_),
    .C(_1394_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3881_ (.A1(_1324_),
    .A2(_1379_),
    .ZN(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3882_ (.A1(_0767_),
    .A2(_1369_),
    .B(_1396_),
    .C(_1394_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3883_ (.I(_0394_),
    .Z(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3884_ (.I(_1397_),
    .Z(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3885_ (.A1(_0363_),
    .A2(_1398_),
    .Z(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3886_ (.A1(_1796_),
    .A2(_0954_),
    .A3(_1399_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3887_ (.I(_1397_),
    .Z(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3888_ (.A1(_0385_),
    .A2(_0391_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3889_ (.A1(_1401_),
    .A2(_0394_),
    .ZN(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3890_ (.I(_1402_),
    .Z(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3891_ (.I(_1403_),
    .Z(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3892_ (.I(_0367_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3893_ (.A1(_0360_),
    .A2(_1400_),
    .B1(_1404_),
    .B2(_1405_),
    .ZN(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3894_ (.A1(_1785_),
    .A2(_1406_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3895_ (.I(_1781_),
    .Z(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3896_ (.A1(_2061_),
    .A2(_1400_),
    .B1(_1404_),
    .B2(_0387_),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3897_ (.A1(_1407_),
    .A2(_1408_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3898_ (.I(_0362_),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3899_ (.A1(\t0pre_counter[3] ),
    .A2(_1400_),
    .B1(_1404_),
    .B2(_1409_),
    .ZN(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3900_ (.A1(_1407_),
    .A2(_1410_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3901_ (.I(_0344_),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3902_ (.A1(_0336_),
    .A2(_1400_),
    .B1(_1404_),
    .B2(_1411_),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3903_ (.A1(_1407_),
    .A2(_1412_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3904_ (.I(_1397_),
    .Z(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3905_ (.I(_1402_),
    .Z(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3906_ (.A1(_0335_),
    .A2(_1413_),
    .B1(_1414_),
    .B2(_0355_),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3907_ (.A1(_1407_),
    .A2(_1415_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3908_ (.I(_1780_),
    .Z(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3909_ (.I(_1416_),
    .Z(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3910_ (.A1(_0334_),
    .A2(_1413_),
    .B1(_1414_),
    .B2(_0349_),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3911_ (.A1(_1417_),
    .A2(_1418_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3912_ (.A1(\t0pre_counter[7] ),
    .A2(_1413_),
    .B1(_1414_),
    .B2(_0340_),
    .ZN(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3913_ (.A1(_1417_),
    .A2(_1419_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3914_ (.I(_0328_),
    .ZN(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3915_ (.A1(_2070_),
    .A2(_1413_),
    .B1(_1414_),
    .B2(_1420_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3916_ (.A1(_1417_),
    .A2(_1421_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3917_ (.I(_1397_),
    .Z(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3918_ (.I(_1402_),
    .Z(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3919_ (.I(_0320_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3920_ (.A1(_2075_),
    .A2(_1422_),
    .B1(_1423_),
    .B2(_1424_),
    .ZN(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3921_ (.A1(_1417_),
    .A2(_1425_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3922_ (.I(_1416_),
    .Z(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3923_ (.I(_2101_),
    .ZN(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3924_ (.A1(_2074_),
    .A2(_1422_),
    .B1(_1423_),
    .B2(_1427_),
    .ZN(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3925_ (.A1(_1426_),
    .A2(_1428_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3926_ (.A1(\t0pre_counter[11] ),
    .A2(_1422_),
    .B1(_1423_),
    .B2(_2099_),
    .ZN(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3927_ (.A1(_1426_),
    .A2(_1429_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3928_ (.A1(_2059_),
    .A2(_1422_),
    .B1(_1423_),
    .B2(_0380_),
    .ZN(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3929_ (.A1(_1426_),
    .A2(_1430_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3930_ (.A1(\t0pre_counter[13] ),
    .A2(_1398_),
    .B1(_1403_),
    .B2(_2084_),
    .ZN(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3931_ (.A1(_1426_),
    .A2(_1431_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3932_ (.I(_1416_),
    .Z(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3933_ (.A1(\t0pre_counter[14] ),
    .A2(_1398_),
    .B1(_1403_),
    .B2(_2068_),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3934_ (.A1(_1432_),
    .A2(_1433_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3935_ (.A1(\t0pre_counter[15] ),
    .A2(_1398_),
    .B1(_1403_),
    .B2(_2078_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3936_ (.A1(_1432_),
    .A2(_1434_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3937_ (.I(_1074_),
    .Z(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3938_ (.A1(_0556_),
    .A2(_1435_),
    .Z(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3939_ (.A1(_1796_),
    .A2(_1071_),
    .A3(_1436_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3940_ (.I(_1435_),
    .Z(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3941_ (.I(_1128_),
    .Z(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3942_ (.I(_0473_),
    .Z(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3943_ (.I(_1439_),
    .Z(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3944_ (.A1(_1440_),
    .A2(_0554_),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3945_ (.A1(_0547_),
    .A2(_1437_),
    .B1(_1438_),
    .B2(_1441_),
    .ZN(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3946_ (.A1(_1432_),
    .A2(_1442_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3947_ (.I(_1439_),
    .Z(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3948_ (.A1(_1443_),
    .A2(_0552_),
    .ZN(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3949_ (.A1(_0476_),
    .A2(_1437_),
    .B1(_1438_),
    .B2(_1444_),
    .ZN(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3950_ (.A1(_1432_),
    .A2(_1445_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3951_ (.I(_1416_),
    .Z(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3952_ (.A1(_1443_),
    .A2(_0550_),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3953_ (.A1(\t1pre_counter[3] ),
    .A2(_1437_),
    .B1(_1438_),
    .B2(_1447_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3954_ (.A1(_1446_),
    .A2(_1448_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3955_ (.A1(_1443_),
    .A2(_0531_),
    .ZN(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3956_ (.A1(_0525_),
    .A2(_1437_),
    .B1(_1438_),
    .B2(_1449_),
    .ZN(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3957_ (.A1(_1446_),
    .A2(_1450_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3958_ (.I(_1435_),
    .Z(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3959_ (.I(_1128_),
    .Z(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3960_ (.A1(_1443_),
    .A2(_0530_),
    .ZN(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3961_ (.A1(_0524_),
    .A2(_1451_),
    .B1(_1452_),
    .B2(_1453_),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3962_ (.A1(_1446_),
    .A2(_1454_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3963_ (.I(_1439_),
    .Z(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3964_ (.A1(_1455_),
    .A2(_0535_),
    .ZN(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3965_ (.A1(_0523_),
    .A2(_1451_),
    .B1(_1452_),
    .B2(_1456_),
    .ZN(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3966_ (.A1(_1446_),
    .A2(_1457_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3967_ (.I(_1784_),
    .Z(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3968_ (.A1(_1455_),
    .A2(_0527_),
    .ZN(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3969_ (.A1(\t1pre_counter[7] ),
    .A2(_1451_),
    .B1(_1452_),
    .B2(_1459_),
    .ZN(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3970_ (.A1(_1458_),
    .A2(_1460_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3971_ (.A1(_1455_),
    .A2(_0519_),
    .ZN(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3972_ (.A1(_0498_),
    .A2(_1451_),
    .B1(_1452_),
    .B2(_1461_),
    .ZN(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3973_ (.A1(_1458_),
    .A2(_1462_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3974_ (.I(_1435_),
    .Z(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3975_ (.I(_1128_),
    .Z(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3976_ (.A1(_1455_),
    .A2(_0510_),
    .ZN(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3977_ (.A1(_0508_),
    .A2(_1463_),
    .B1(_1464_),
    .B2(_1465_),
    .ZN(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3978_ (.A1(_1458_),
    .A2(_1466_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3979_ (.I(_1439_),
    .Z(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3980_ (.A1(_1467_),
    .A2(_0502_),
    .ZN(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3981_ (.A1(_0497_),
    .A2(_1463_),
    .B1(_1464_),
    .B2(_1468_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3982_ (.A1(_1458_),
    .A2(_1469_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3983_ (.I(_1784_),
    .Z(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3984_ (.A1(_1467_),
    .A2(_0569_),
    .ZN(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3985_ (.A1(\t1pre_counter[11] ),
    .A2(_1463_),
    .B1(_1464_),
    .B2(_1471_),
    .ZN(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3986_ (.A1(_1470_),
    .A2(_1472_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3987_ (.A1(_1467_),
    .A2(_0564_),
    .ZN(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3988_ (.A1(\t1pre_counter[12] ),
    .A2(_1463_),
    .B1(_1464_),
    .B2(_1473_),
    .ZN(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3989_ (.A1(_1470_),
    .A2(_1474_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3990_ (.A1(_1467_),
    .A2(_0489_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3991_ (.A1(\t1pre_counter[13] ),
    .A2(_1440_),
    .B1(_1077_),
    .B2(_1475_),
    .ZN(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3992_ (.A1(_1470_),
    .A2(_1476_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3993_ (.A1(_1075_),
    .A2(_0481_),
    .ZN(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3994_ (.A1(\t1pre_counter[14] ),
    .A2(_1440_),
    .B1(_1077_),
    .B2(_1477_),
    .ZN(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3995_ (.A1(_1470_),
    .A2(_1478_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3996_ (.A1(_1075_),
    .A2(_0483_),
    .ZN(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3997_ (.A1(\t1pre_counter[15] ),
    .A2(_1440_),
    .B1(_1077_),
    .B2(_1479_),
    .ZN(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3998_ (.A1(_0740_),
    .A2(_1480_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3999_ (.A1(_1890_),
    .A2(_1854_),
    .A3(_0459_),
    .ZN(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4000_ (.I(_1481_),
    .Z(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4001_ (.I(_1482_),
    .Z(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4002_ (.A1(_1056_),
    .A2(_1483_),
    .ZN(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4003_ (.A1(_0855_),
    .A2(_0862_),
    .ZN(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4004_ (.A1(_1485_),
    .A2(_0941_),
    .ZN(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4005_ (.I(_1486_),
    .Z(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4006_ (.A1(_0855_),
    .A2(_0862_),
    .Z(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4007_ (.I(_1488_),
    .Z(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4008_ (.A1(_1239_),
    .A2(_1489_),
    .ZN(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4009_ (.A1(_1892_),
    .A2(_1273_),
    .ZN(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4010_ (.A1(_1239_),
    .A2(_1487_),
    .B(_1490_),
    .C(_1491_),
    .ZN(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4011_ (.A1(_1484_),
    .A2(_1492_),
    .B(_1371_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4012_ (.I(_1481_),
    .Z(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4013_ (.I(_1493_),
    .Z(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4014_ (.A1(_1243_),
    .A2(_0943_),
    .A3(_1490_),
    .ZN(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4015_ (.I(_1486_),
    .Z(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4016_ (.A1(_1243_),
    .A2(_1240_),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4017_ (.I(_1482_),
    .Z(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4018_ (.A1(_1496_),
    .A2(_1497_),
    .B(_1498_),
    .ZN(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4019_ (.A1(_1283_),
    .A2(_1494_),
    .B1(_1495_),
    .B2(_1499_),
    .C(_1161_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4020_ (.I(_1482_),
    .Z(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4021_ (.I(_1500_),
    .Z(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4022_ (.I(_1485_),
    .Z(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4023_ (.A1(_0908_),
    .A2(_0911_),
    .ZN(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4024_ (.I(_0942_),
    .Z(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4025_ (.A1(_1502_),
    .A2(_1503_),
    .B(_1504_),
    .C(_0935_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4026_ (.A1(_0935_),
    .A2(_1503_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4027_ (.A1(_1496_),
    .A2(_1506_),
    .B(_1498_),
    .ZN(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4028_ (.A1(_1290_),
    .A2(_1501_),
    .B1(_1505_),
    .B2(_1507_),
    .C(_1161_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4029_ (.A1(_0935_),
    .A2(_1243_),
    .A3(_1239_),
    .A4(_1489_),
    .ZN(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4030_ (.A1(_0902_),
    .A2(_0943_),
    .A3(_1508_),
    .ZN(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4031_ (.I(_1486_),
    .Z(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4032_ (.A1(_0902_),
    .A2(_0906_),
    .A3(_1503_),
    .ZN(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4033_ (.A1(_1510_),
    .A2(_1511_),
    .B(_1498_),
    .ZN(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4034_ (.A1(_0979_),
    .A2(_1501_),
    .B1(_1509_),
    .B2(_1512_),
    .C(_1161_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4035_ (.I(_0941_),
    .Z(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4036_ (.I(_1513_),
    .Z(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4037_ (.A1(\timer2[3] ),
    .A2(\timer2[2] ),
    .A3(_0908_),
    .A4(\timer2[0] ),
    .Z(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4038_ (.I(_1488_),
    .Z(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4039_ (.I(_1516_),
    .Z(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4040_ (.A1(_1514_),
    .A2(_1515_),
    .B(_1517_),
    .ZN(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4041_ (.A1(_0915_),
    .A2(_1515_),
    .Z(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4042_ (.A1(\timer2[4] ),
    .A2(_1518_),
    .B1(_1519_),
    .B2(_1487_),
    .C(_1483_),
    .ZN(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4043_ (.I(_1491_),
    .Z(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4044_ (.I(_1804_),
    .Z(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4045_ (.A1(_1296_),
    .A2(_1521_),
    .B(_1522_),
    .ZN(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4046_ (.A1(_1520_),
    .A2(_1523_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4047_ (.A1(\timer2[4] ),
    .A2(_1515_),
    .Z(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4048_ (.I(_1524_),
    .Z(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4049_ (.A1(_1513_),
    .A2(_1525_),
    .B(_1516_),
    .ZN(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4050_ (.A1(_0919_),
    .A2(_1525_),
    .Z(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4051_ (.I(_1486_),
    .Z(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4052_ (.A1(_0898_),
    .A2(_1526_),
    .B1(_1527_),
    .B2(_1528_),
    .C(_1493_),
    .ZN(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4053_ (.I(_0987_),
    .Z(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4054_ (.A1(_1299_),
    .A2(_1494_),
    .B(_1529_),
    .C(_1530_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4055_ (.A1(_0898_),
    .A2(_1525_),
    .ZN(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4056_ (.A1(_1502_),
    .A2(_1531_),
    .B(_1504_),
    .C(_0893_),
    .ZN(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4057_ (.A1(_0893_),
    .A2(_1531_),
    .ZN(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4058_ (.A1(_1510_),
    .A2(_1533_),
    .B(_1498_),
    .ZN(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4059_ (.I(_1006_),
    .Z(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4060_ (.A1(_1001_),
    .A2(_1501_),
    .B1(_1532_),
    .B2(_1534_),
    .C(_1535_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4061_ (.A1(_0893_),
    .A2(_0898_),
    .A3(_1489_),
    .A4(_1525_),
    .ZN(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4062_ (.A1(_0892_),
    .A2(_1504_),
    .A3(_1536_),
    .ZN(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4063_ (.A1(_0892_),
    .A2(_0921_),
    .A3(_1531_),
    .ZN(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4064_ (.A1(_1510_),
    .A2(_1538_),
    .B(_1500_),
    .ZN(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4065_ (.A1(_1305_),
    .A2(_1501_),
    .B1(_1537_),
    .B2(_1539_),
    .C(_1535_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4066_ (.A1(_0892_),
    .A2(\timer2[6] ),
    .A3(\timer2[5] ),
    .A4(_1524_),
    .Z(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4067_ (.A1(_1514_),
    .A2(_1540_),
    .B(_1517_),
    .ZN(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4068_ (.I(_1540_),
    .ZN(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4069_ (.A1(_0874_),
    .A2(_1542_),
    .ZN(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4070_ (.I(_1482_),
    .Z(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4071_ (.A1(_0874_),
    .A2(_1541_),
    .B1(_1543_),
    .B2(_1487_),
    .C(_1544_),
    .ZN(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4072_ (.I(_0723_),
    .Z(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4073_ (.A1(_1546_),
    .A2(_1521_),
    .B(_1522_),
    .ZN(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4074_ (.A1(_1545_),
    .A2(_1547_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4075_ (.A1(_0874_),
    .A2(_1540_),
    .Z(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4076_ (.A1(_1513_),
    .A2(_1548_),
    .B(_1516_),
    .ZN(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4077_ (.A1(_1261_),
    .A2(_0930_),
    .A3(_1542_),
    .ZN(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4078_ (.A1(_1261_),
    .A2(_1549_),
    .B1(_1550_),
    .B2(_1528_),
    .C(_1493_),
    .ZN(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4079_ (.A1(_1020_),
    .A2(_1494_),
    .B(_1551_),
    .C(_1530_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4080_ (.A1(_1261_),
    .A2(_1548_),
    .ZN(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4081_ (.A1(_1502_),
    .A2(_1552_),
    .B(_1504_),
    .C(_1264_),
    .ZN(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4082_ (.A1(_1264_),
    .A2(_1552_),
    .ZN(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4083_ (.A1(_1510_),
    .A2(_1554_),
    .B(_1500_),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4084_ (.A1(_1023_),
    .A2(_1483_),
    .B1(_1553_),
    .B2(_1555_),
    .C(_1535_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4085_ (.A1(_1264_),
    .A2(_0873_),
    .A3(_1548_),
    .Z(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4086_ (.A1(_1514_),
    .A2(_1556_),
    .B(_1517_),
    .ZN(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4087_ (.A1(_0870_),
    .A2(_1556_),
    .Z(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4088_ (.A1(\timer2[11] ),
    .A2(_1557_),
    .B1(_1558_),
    .B2(_1487_),
    .C(_1544_),
    .ZN(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4089_ (.A1(_1354_),
    .A2(_1521_),
    .B(_1522_),
    .ZN(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4090_ (.A1(_1559_),
    .A2(_1560_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4091_ (.A1(\timer2[11] ),
    .A2(\timer2[10] ),
    .A3(_0873_),
    .A4(_1548_),
    .Z(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4092_ (.A1(_1514_),
    .A2(_1561_),
    .B(_1489_),
    .ZN(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4093_ (.A1(_0883_),
    .A2(_1561_),
    .Z(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4094_ (.A1(\timer2[12] ),
    .A2(_1562_),
    .B1(_1563_),
    .B2(_1496_),
    .C(_1544_),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4095_ (.A1(_1315_),
    .A2(_1521_),
    .B(_1522_),
    .ZN(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4096_ (.A1(_1564_),
    .A2(_1565_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4097_ (.A1(\timer2[12] ),
    .A2(_1561_),
    .ZN(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4098_ (.A1(_1485_),
    .A2(_1566_),
    .B(_0942_),
    .C(\timer2[13] ),
    .ZN(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4099_ (.A1(\timer2[13] ),
    .A2(_1566_),
    .ZN(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4100_ (.A1(_1528_),
    .A2(_1568_),
    .B(_1500_),
    .ZN(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4101_ (.A1(_1041_),
    .A2(_1483_),
    .B1(_1567_),
    .B2(_1569_),
    .C(_1535_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4102_ (.A1(_0882_),
    .A2(_1566_),
    .ZN(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4103_ (.A1(_1513_),
    .A2(_1570_),
    .B(_1516_),
    .ZN(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4104_ (.I(_1570_),
    .ZN(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4105_ (.A1(_0886_),
    .A2(_1572_),
    .ZN(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4106_ (.A1(_0886_),
    .A2(_1571_),
    .B1(_1573_),
    .B2(_1528_),
    .C(_1493_),
    .ZN(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4107_ (.A1(_1046_),
    .A2(_1494_),
    .B(_1574_),
    .C(_1530_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4108_ (.A1(_0886_),
    .A2(_1517_),
    .A3(_1570_),
    .ZN(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4109_ (.A1(_0864_),
    .A2(_0942_),
    .Z(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4110_ (.A1(_0864_),
    .A2(_0865_),
    .A3(_1572_),
    .ZN(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4111_ (.A1(_1575_),
    .A2(_1576_),
    .B1(_1577_),
    .B2(_1496_),
    .C(_1544_),
    .ZN(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4112_ (.A1(_1324_),
    .A2(_1491_),
    .B(_1805_),
    .ZN(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4113_ (.A1(_1578_),
    .A2(_1579_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4114_ (.A1(_1862_),
    .A2(_1273_),
    .ZN(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4115_ (.I(_1580_),
    .Z(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4116_ (.A1(\t0_top[0] ),
    .A2(_1581_),
    .ZN(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4117_ (.A1(_1869_),
    .A2(_1884_),
    .A3(_1278_),
    .ZN(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4118_ (.I(_1583_),
    .Z(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4119_ (.I(_1584_),
    .Z(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4120_ (.A1(_1277_),
    .A2(_1585_),
    .ZN(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4121_ (.A1(_0646_),
    .A2(_1582_),
    .A3(_1586_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4122_ (.I(_1580_),
    .Z(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4123_ (.A1(\t0_top[1] ),
    .A2(_1581_),
    .ZN(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4124_ (.A1(_1284_),
    .A2(_1587_),
    .B(_1588_),
    .C(_1394_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4125_ (.I(_1583_),
    .Z(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4126_ (.I(_1589_),
    .Z(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4127_ (.I(_1584_),
    .Z(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4128_ (.A1(_0976_),
    .A2(_1591_),
    .ZN(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4129_ (.I(_1317_),
    .Z(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4130_ (.I(_1593_),
    .Z(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4131_ (.A1(_0407_),
    .A2(_1590_),
    .B(_1592_),
    .C(_1594_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4132_ (.A1(\t0_top[3] ),
    .A2(_1581_),
    .ZN(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4133_ (.A1(_1292_),
    .A2(_1587_),
    .B(_1595_),
    .C(_1594_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4134_ (.A1(_0989_),
    .A2(_1591_),
    .ZN(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4135_ (.A1(_0404_),
    .A2(_1590_),
    .B(_1596_),
    .C(_1594_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4136_ (.A1(\temp[5] ),
    .A2(_1591_),
    .ZN(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4137_ (.A1(_0403_),
    .A2(_1590_),
    .B(_1597_),
    .C(_1594_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4138_ (.A1(\temp[6] ),
    .A2(_1591_),
    .ZN(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4139_ (.I(_1593_),
    .Z(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4140_ (.A1(_0400_),
    .A2(_1590_),
    .B(_1598_),
    .C(_1599_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4141_ (.I(_1584_),
    .Z(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4142_ (.I(_1584_),
    .Z(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4143_ (.A1(_1008_),
    .A2(_1601_),
    .ZN(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4144_ (.A1(_0397_),
    .A2(_1600_),
    .B(_1602_),
    .C(_1599_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4145_ (.A1(_1546_),
    .A2(_1601_),
    .ZN(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4146_ (.A1(_0430_),
    .A2(_1600_),
    .B(_1603_),
    .C(_1599_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4147_ (.I(_0728_),
    .Z(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4148_ (.A1(\t0_top[9] ),
    .A2(_1581_),
    .ZN(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4149_ (.A1(_1604_),
    .A2(_1587_),
    .B(_1605_),
    .C(_1599_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4150_ (.A1(net11),
    .A2(_1601_),
    .ZN(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4151_ (.I(_1593_),
    .Z(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4152_ (.A1(_0421_),
    .A2(_1600_),
    .B(_1606_),
    .C(_1607_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4153_ (.A1(_1028_),
    .A2(_1601_),
    .ZN(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4154_ (.A1(_0419_),
    .A2(_1600_),
    .B(_1608_),
    .C(_1607_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4155_ (.A1(_0469_),
    .A2(_1589_),
    .ZN(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4156_ (.A1(_0444_),
    .A2(_1585_),
    .B(_1609_),
    .C(_1607_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4157_ (.I(_0944_),
    .Z(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4158_ (.A1(\t0_top[13] ),
    .A2(_1580_),
    .ZN(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4159_ (.A1(_1610_),
    .A2(_1587_),
    .B(_1611_),
    .C(_1607_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4160_ (.A1(_1322_),
    .A2(_1589_),
    .ZN(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4161_ (.I(_1593_),
    .Z(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4162_ (.A1(_0440_),
    .A2(_1585_),
    .B(_1612_),
    .C(_1613_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4163_ (.I(_0738_),
    .Z(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4164_ (.A1(_1614_),
    .A2(_1589_),
    .ZN(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4165_ (.A1(_0438_),
    .A2(_1585_),
    .B(_1615_),
    .C(_1613_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4166_ (.A1(_0949_),
    .A2(_1884_),
    .A3(_0460_),
    .ZN(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4167_ (.I(_1616_),
    .Z(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4168_ (.I(_1617_),
    .Z(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4169_ (.I(_1617_),
    .Z(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4170_ (.A1(_1056_),
    .A2(_1619_),
    .ZN(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4171_ (.A1(_0618_),
    .A2(_1618_),
    .B(_1620_),
    .C(_1613_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4172_ (.I(_1616_),
    .Z(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4173_ (.A1(_0962_),
    .A2(_1621_),
    .ZN(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4174_ (.A1(_0616_),
    .A2(_1618_),
    .B(_1622_),
    .C(_1613_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4175_ (.A1(_1903_),
    .A2(_0719_),
    .ZN(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4176_ (.I(_1623_),
    .Z(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4177_ (.A1(\t1_top[2] ),
    .A2(_1624_),
    .ZN(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4178_ (.A1(_0976_),
    .A2(_1619_),
    .ZN(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4179_ (.A1(_0646_),
    .A2(_1625_),
    .A3(_1626_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4180_ (.I(_1623_),
    .Z(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4181_ (.I(_1627_),
    .Z(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4182_ (.A1(\t1_top[3] ),
    .A2(_1624_),
    .ZN(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4183_ (.I(_0464_),
    .Z(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4184_ (.I(_1630_),
    .Z(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4185_ (.A1(_0980_),
    .A2(_1628_),
    .B(_1629_),
    .C(_1631_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4186_ (.A1(_0989_),
    .A2(_1621_),
    .ZN(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4187_ (.A1(_0613_),
    .A2(_1618_),
    .B(_1632_),
    .C(_1631_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4188_ (.A1(\temp[5] ),
    .A2(_1621_),
    .ZN(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4189_ (.A1(_0625_),
    .A2(_1618_),
    .B(_1633_),
    .C(_1631_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4190_ (.A1(\t1_top[6] ),
    .A2(_1624_),
    .ZN(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4191_ (.A1(_1301_),
    .A2(_1628_),
    .B(_1634_),
    .C(_1631_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4192_ (.A1(\t1_top[7] ),
    .A2(_1627_),
    .ZN(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4193_ (.I(_1630_),
    .Z(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4194_ (.A1(_1306_),
    .A2(_1628_),
    .B(_1635_),
    .C(_1636_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4195_ (.I(\t1_top[8] ),
    .ZN(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4196_ (.I(_1617_),
    .Z(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4197_ (.A1(_1308_),
    .A2(_1621_),
    .ZN(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4198_ (.A1(_1637_),
    .A2(_1638_),
    .B(_1639_),
    .C(_1636_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4199_ (.A1(\t1_top[9] ),
    .A2(_1627_),
    .ZN(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4200_ (.A1(_1020_),
    .A2(_1628_),
    .B(_1640_),
    .C(_1636_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4201_ (.A1(\t1_top[10] ),
    .A2(_1627_),
    .ZN(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4202_ (.A1(_1023_),
    .A2(_1624_),
    .B(_1641_),
    .C(_1636_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4203_ (.I(_1616_),
    .Z(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4204_ (.A1(_1028_),
    .A2(_1642_),
    .ZN(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4205_ (.I(_1630_),
    .Z(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4206_ (.A1(_0593_),
    .A2(_1638_),
    .B(_1643_),
    .C(_1644_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4207_ (.A1(_0469_),
    .A2(_1642_),
    .ZN(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4208_ (.D(_0000_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\pwm_ctr2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4209_ (.D(_0001_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\pwm_ctr2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4210_ (.D(_0002_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\pwm_ctr2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4211_ (.D(_0003_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\pwm_ctr2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4212_ (.D(_0004_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\pwm_ctr2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4213_ (.D(_0005_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\pwm_ctr2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4214_ (.D(_0006_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\pwm_ctr2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4215_ (.D(_0007_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\pwm_ctr2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4216_ (.D(_0008_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4217_ (.D(_0009_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4218_ (.D(_0010_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4219_ (.D(_0011_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4220_ (.D(_0012_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4221_ (.D(_0013_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4222_ (.D(_0014_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4223_ (.D(_0015_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4224_ (.D(_0016_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4225_ (.D(_0017_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4226_ (.D(_0018_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(net34));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4227_ (.D(_0019_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(net35));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4228_ (.D(_0020_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4229_ (.D(_0021_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4230_ (.D(_0022_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4231_ (.D(_0023_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\settings[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4232_ (.D(_0024_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\settings[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4233_ (.D(_0025_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\settings[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4234_ (.D(_0026_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(tmr0_ext));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4235_ (.D(_0027_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(tmr1_ext));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4236_ (.D(_0028_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4237_ (.D(_0029_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(last_tmr0_clk));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4238_ (.D(_0030_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(last_tmr1_clk));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4239_ (.D(_0031_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\timer0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4240_ (.D(_0032_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\timer0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4241_ (.D(_0033_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\timer0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4242_ (.D(_0034_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\timer0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4243_ (.D(_0035_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\timer0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4244_ (.D(_0036_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\timer0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4245_ (.D(_0037_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\timer0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4246_ (.D(_0038_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\timer0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4247_ (.D(_0039_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\timer0[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4248_ (.D(_0040_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\timer0[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4249_ (.D(_0041_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\timer0[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4250_ (.D(_0042_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\timer0[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4251_ (.D(_0043_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\timer0[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4252_ (.D(_0044_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\timer0[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4253_ (.D(_0045_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\timer0[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4254_ (.D(_0046_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\timer0[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4255_ (.D(_0047_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\timer1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4256_ (.D(_0048_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\timer1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4257_ (.D(_0049_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\timer1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4258_ (.D(_0050_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\timer1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4259_ (.D(_0051_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\timer1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4260_ (.D(_0052_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\timer1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4261_ (.D(_0053_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\timer1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4262_ (.D(_0054_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\timer1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4263_ (.D(_0055_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\timer1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4264_ (.D(_0056_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\timer1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4265_ (.D(_0057_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\timer1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4266_ (.D(_0058_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\timer1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4267_ (.D(_0059_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\timer1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4268_ (.D(_0060_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\timer1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4269_ (.D(_0061_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\timer1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4270_ (.D(_0062_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\timer1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4271_ (.D(_0063_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\t0_capture[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4272_ (.D(_0064_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\t0_capture[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4273_ (.D(_0065_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\t0_capture[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4274_ (.D(_0066_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\t0_capture[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4275_ (.D(_0067_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\t0_capture[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4276_ (.D(_0068_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\t0_capture[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4277_ (.D(_0069_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\t0_capture[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4278_ (.D(_0070_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\t0_capture[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4279_ (.D(_0071_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\t0_capture[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4280_ (.D(_0072_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\t0_capture[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4281_ (.D(_0073_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\t0_capture[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4282_ (.D(_0074_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\t0_capture[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4283_ (.D(_0075_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\t0_capture[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4284_ (.D(_0076_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\t0_capture[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4285_ (.D(_0077_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\t0_capture[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4286_ (.D(_0078_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\t0_capture[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4287_ (.D(_0079_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\t1_capture[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4288_ (.D(_0080_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\t1_capture[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4289_ (.D(_0081_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\t1_capture[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4290_ (.D(_0082_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\t1_capture[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4291_ (.D(_0083_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\t1_capture[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4292_ (.D(_0084_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\t1_capture[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4293_ (.D(_0085_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\t1_capture[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4294_ (.D(_0086_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\t1_capture[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4295_ (.D(_0087_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\t1_capture[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4296_ (.D(_0088_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\t1_capture[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4297_ (.D(_0089_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\t1_capture[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4298_ (.D(_0090_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\t1_capture[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4299_ (.D(_0091_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\t1_capture[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4300_ (.D(_0092_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\t1_capture[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4301_ (.D(_0093_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\t1_capture[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4302_ (.D(_0094_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\t1_capture[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4303_ (.D(_0095_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\t2_capture[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4304_ (.D(_0096_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\t2_capture[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4305_ (.D(_0097_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\t2_capture[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4306_ (.D(_0098_),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(\t2_capture[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4307_ (.D(_0099_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\t2_capture[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4308_ (.D(_0100_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\t2_capture[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4309_ (.D(_0101_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\t2_capture[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4310_ (.D(_0102_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\t2_capture[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4311_ (.D(_0103_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\t2_capture[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4312_ (.D(_0104_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\t2_capture[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4313_ (.D(_0105_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\t2_capture[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4314_ (.D(_0106_),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(\t2_capture[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4315_ (.D(_0107_),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(\t2_capture[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4316_ (.D(_0108_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\t2_capture[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4317_ (.D(_0109_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\t2_capture[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4318_ (.D(_0110_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\t2_capture[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4319_ (.D(_0111_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\t0pre[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4320_ (.D(_0112_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\t0pre[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4321_ (.D(_0113_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\t0pre[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4322_ (.D(_0114_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\t0pre[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4323_ (.D(_0115_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\t0pre[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4324_ (.D(_0116_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\t0pre[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4325_ (.D(_0117_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\t0pre[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4326_ (.D(_0118_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\t0pre[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4327_ (.D(_0119_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\t0pre[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4328_ (.D(_0120_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\t0pre[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4329_ (.D(_0121_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\t0pre[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4330_ (.D(_0122_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\t0pre[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4331_ (.D(_0123_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\t0pre[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4332_ (.D(_0124_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\t0pre[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4333_ (.D(_0125_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\t0pre[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4334_ (.D(_0126_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\t0pre[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4335_ (.D(_0127_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\t1pre[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4336_ (.D(_0128_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\t1pre[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4337_ (.D(_0129_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\t1pre[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4338_ (.D(_0130_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\t1pre[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4339_ (.D(_0131_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\t1pre[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4340_ (.D(_0132_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\t1pre[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4341_ (.D(_0133_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\t1pre[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4342_ (.D(_0134_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\t1pre[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4343_ (.D(_0135_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\t1pre[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4344_ (.D(_0136_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\t1pre[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4345_ (.D(_0137_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\t1pre[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4346_ (.D(_0138_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\t1pre[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4347_ (.D(_0139_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\t1pre[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4348_ (.D(_0140_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\t1pre[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4349_ (.D(_0141_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\t1pre[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4350_ (.D(_0142_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\t1pre[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4351_ (.D(_0143_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\t2pre[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4352_ (.D(_0144_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\t2pre[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4353_ (.D(_0145_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\t2pre[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4354_ (.D(_0146_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\t2pre[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4355_ (.D(_0147_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\t2pre[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4356_ (.D(_0148_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\t2pre[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4357_ (.D(_0149_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\t2pre[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4358_ (.D(_0150_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\t2pre[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4359_ (.D(_0151_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\t2pre[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4360_ (.D(_0152_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\t2pre[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4361_ (.D(_0153_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\t2pre[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4362_ (.D(_0154_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\t2pre[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4363_ (.D(_0155_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\t2pre[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4364_ (.D(_0156_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\t2pre[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4365_ (.D(_0157_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\t2pre[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4366_ (.D(_0158_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\t2pre[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4367_ (.D(_0159_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\t0pre_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4368_ (.D(_0160_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\t0pre_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4369_ (.D(_0161_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\t0pre_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4370_ (.D(_0162_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\t0pre_counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4371_ (.D(_0163_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\t0pre_counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4372_ (.D(_0164_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\t0pre_counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4373_ (.D(_0165_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\t0pre_counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4374_ (.D(_0166_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\t0pre_counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4375_ (.D(_0167_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\t0pre_counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4376_ (.D(_0168_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\t0pre_counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4377_ (.D(_0169_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\t0pre_counter[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4378_ (.D(_0170_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\t0pre_counter[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4379_ (.D(_0171_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\t0pre_counter[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4380_ (.D(_0172_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\t0pre_counter[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4381_ (.D(_0173_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\t0pre_counter[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4382_ (.D(_0174_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\t0pre_counter[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4383_ (.D(_0175_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\t1pre_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4384_ (.D(_0176_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\t1pre_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4385_ (.D(_0177_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\t1pre_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4386_ (.D(_0178_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\t1pre_counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4387_ (.D(_0179_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\t1pre_counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4388_ (.D(_0180_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\t1pre_counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4389_ (.D(_0181_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\t1pre_counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4390_ (.D(_0182_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\t1pre_counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4391_ (.D(_0183_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\t1pre_counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4392_ (.D(_0184_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\t1pre_counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4393_ (.D(_0185_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\t1pre_counter[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4394_ (.D(_0186_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\t1pre_counter[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4395_ (.D(_0187_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\t1pre_counter[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4396_ (.D(_0188_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\t1pre_counter[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4397_ (.D(_0189_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\t1pre_counter[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4398_ (.D(_0190_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\t1pre_counter[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4399_ (.D(_0191_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\timer2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4400_ (.D(_0192_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\timer2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4401_ (.D(_0193_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\timer2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4402_ (.D(_0194_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\timer2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4403_ (.D(_0195_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\timer2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4404_ (.D(_0196_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\timer2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4405_ (.D(_0197_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\timer2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4406_ (.D(_0198_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\timer2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4407_ (.D(_0199_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\timer2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4408_ (.D(_0200_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\timer2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4409_ (.D(_0201_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\timer2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4410_ (.D(_0202_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\timer2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4411_ (.D(_0203_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\timer2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4412_ (.D(_0204_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(\timer2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4413_ (.D(_0205_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\timer2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4414_ (.D(_0206_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\timer2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4415_ (.D(_0207_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\t0_top[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4416_ (.D(_0208_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\t0_top[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4417_ (.D(_0209_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\t0_top[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4418_ (.D(_0210_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\t0_top[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4419_ (.D(_0211_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\t0_top[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4420_ (.D(_0212_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\t0_top[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4421_ (.D(_0213_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\t0_top[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4422_ (.D(_0214_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\t0_top[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4423_ (.D(_0215_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\t0_top[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4424_ (.D(_0216_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\t0_top[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4425_ (.D(_0217_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\t0_top[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4426_ (.D(_0218_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\t0_top[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4427_ (.D(_0219_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\t0_top[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4428_ (.D(_0220_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\t0_top[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4429_ (.D(_0221_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\t0_top[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4430_ (.D(_0222_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\t0_top[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4431_ (.D(_0223_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\t1_top[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4432_ (.D(_0224_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\t1_top[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4433_ (.D(_0225_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\t1_top[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4434_ (.D(_0226_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\t1_top[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4435_ (.D(_0227_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\t1_top[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4436_ (.D(_0228_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\t1_top[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4437_ (.D(_0229_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\t1_top[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4438_ (.D(_0230_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\t1_top[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4439_ (.D(_0231_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\t1_top[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4440_ (.D(_0232_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\t1_top[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4441_ (.D(_0233_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\t1_top[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4442_ (.D(_0234_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\t1_top[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4443_ (.D(_0235_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\t1_top[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4444_ (.D(_0236_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\t1_top[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4445_ (.D(_0237_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\t1_top[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4446_ (.D(_0238_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\t1_top[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4447_ (.D(_0239_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\t2_top[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4448_ (.D(_0240_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\t2_top[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4449_ (.D(_0241_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\t2_top[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4450_ (.D(_0242_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\t2_top[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4451_ (.D(_0243_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\t2_top[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4452_ (.D(_0244_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\t2_top[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4453_ (.D(_0245_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(\t2_top[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4454_ (.D(_0246_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\t2_top[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4455_ (.D(_0247_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\t2_top[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4456_ (.D(_0248_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\t2_top[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4457_ (.D(_0249_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\t2_top[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4458_ (.D(_0250_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\t2_top[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4459_ (.D(_0251_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\t2_top[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4460_ (.D(_0252_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\t2_top[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4461_ (.D(_0253_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\t2_top[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4462_ (.D(_0254_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\t2_top[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4463_ (.D(_0255_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\t2pre_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4464_ (.D(_0256_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\t2pre_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4465_ (.D(_0257_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\t2pre_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4466_ (.D(_0258_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\t2pre_counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4467_ (.D(_0259_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\t2pre_counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4468_ (.D(_0260_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\t2pre_counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4469_ (.D(_0261_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\t2pre_counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4470_ (.D(_0262_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\t2pre_counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4471_ (.D(_0263_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\t2pre_counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4472_ (.D(_0264_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\t2pre_counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4473_ (.D(_0265_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\t2pre_counter[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4474_ (.D(_0266_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\t2pre_counter[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4475_ (.D(_0267_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\t2pre_counter[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4476_ (.D(_0268_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\t2pre_counter[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4477_ (.D(_0269_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\t2pre_counter[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4478_ (.D(_0270_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\t2pre_counter[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4479_ (.D(_0271_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\pwm_ctr0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4480_ (.D(_0272_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\pwm_ctr0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4481_ (.D(_0273_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\pwm_ctr0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4482_ (.D(_0274_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\pwm_ctr0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4483_ (.D(_0275_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\pwm_ctr0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4484_ (.D(_0276_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\pwm_ctr0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4485_ (.D(_0277_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\pwm_ctr0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4486_ (.D(_0278_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\pwm_ctr0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4487_ (.D(_0279_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\pwm_ctr1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4488_ (.D(_0280_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\pwm_ctr1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4489_ (.D(_0281_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\pwm_ctr1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4490_ (.D(_0282_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\pwm_ctr1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4491_ (.D(_0283_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\pwm_ctr1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4492_ (.D(_0284_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\pwm_ctr1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4493_ (.D(_0285_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\pwm_ctr1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4494_ (.D(_0286_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\pwm_ctr1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4495_ (.D(_0287_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\pw0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4496_ (.D(_0288_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\pw0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4497_ (.D(_0289_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\pw0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4498_ (.D(_0290_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\pw0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4499_ (.D(_0291_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\pw0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4500_ (.D(_0292_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\pw0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4501_ (.D(_0293_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\pw0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4502_ (.D(_0294_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\pw0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4503_ (.D(_0295_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\pw1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4504_ (.D(_0296_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\pw1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4505_ (.D(_0297_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\pw1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4506_ (.D(_0298_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\pw1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4507_ (.D(_0299_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\pw1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4508_ (.D(_0300_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\pw1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4509_ (.D(_0301_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\pw1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4510_ (.D(_0302_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\pw1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4511_ (.D(_0303_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\pw2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4512_ (.D(_0304_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\pw2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4513_ (.D(_0305_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\pw2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4514_ (.D(_0306_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\pw2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4515_ (.D(_0307_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\pw2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4516_ (.D(_0308_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\pw2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4517_ (.D(_0309_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\pw2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4518_ (.D(_0310_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\pw2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4519_ (.D(_0311_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\temp[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4520_ (.D(_0312_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\temp[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4521_ (.D(_0313_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\temp[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4522_ (.D(_0314_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\temp[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4523_ (.D(_0315_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\temp[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4524_ (.D(_0316_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\temp[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4525_ (.D(_0317_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\temp[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4526_ (.D(_0318_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\temp[7] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_0__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_1__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_2__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_3__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_4__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_5__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_6__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_7__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.I(clknet_3_3__leaf_wb_clk_i),
    .Z(clknet_leaf_10_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.I(clknet_3_3__leaf_wb_clk_i),
    .Z(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.I(clknet_3_3__leaf_wb_clk_i),
    .Z(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.I(clknet_3_2__leaf_wb_clk_i),
    .Z(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.I(clknet_3_2__leaf_wb_clk_i),
    .Z(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.I(clknet_3_3__leaf_wb_clk_i),
    .Z(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.I(clknet_3_2__leaf_wb_clk_i),
    .Z(clknet_leaf_16_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.I(clknet_3_2__leaf_wb_clk_i),
    .Z(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.I(clknet_3_2__leaf_wb_clk_i),
    .Z(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.I(clknet_3_2__leaf_wb_clk_i),
    .Z(clknet_leaf_19_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.I(clknet_3_2__leaf_wb_clk_i),
    .Z(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.I(clknet_3_2__leaf_wb_clk_i),
    .Z(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.I(clknet_3_2__leaf_wb_clk_i),
    .Z(clknet_leaf_22_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.I(clknet_3_2__leaf_wb_clk_i),
    .Z(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.I(clknet_3_2__leaf_wb_clk_i),
    .Z(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.I(clknet_3_3__leaf_wb_clk_i),
    .Z(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.I(clknet_3_3__leaf_wb_clk_i),
    .Z(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.I(clknet_3_3__leaf_wb_clk_i),
    .Z(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.I(clknet_3_3__leaf_wb_clk_i),
    .Z(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.I(clknet_3_3__leaf_wb_clk_i),
    .Z(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.I(clknet_3_3__leaf_wb_clk_i),
    .Z(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.I(clknet_3_3__leaf_wb_clk_i),
    .Z(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.I(clknet_3_3__leaf_wb_clk_i),
    .Z(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_72_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_78_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_81_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_81_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_82_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_82_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_83_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_83_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_84_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_84_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_85_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_85_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_86_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_86_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_87_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_87_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_88_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_88_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_89_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_89_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_8_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_90_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_90_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_91_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_91_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_92_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_92_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_93_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_93_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1 (.I(addr[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input10 (.I(data_in[1]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input11 (.I(data_in[2]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input12 (.I(data_in[3]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input13 (.I(data_in[4]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input14 (.I(data_in[5]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input15 (.I(data_in[6]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(data_in[7]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input17 (.I(rst),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input18 (.I(tmr0_clk),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input19 (.I(tmr1_clk),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input2 (.I(addr[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input3 (.I(addr[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input4 (.I(addr[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input5 (.I(addr[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input6 (.I(addr[5]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input7 (.I(bus_cyc),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input8 (.I(bus_we),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(data_in[0]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output20 (.I(net20),
    .Z(data_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output21 (.I(net21),
    .Z(data_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output22 (.I(net22),
    .Z(data_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output23 (.I(net23),
    .Z(data_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output24 (.I(net24),
    .Z(data_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output25 (.I(net25),
    .Z(data_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output26 (.I(net26),
    .Z(data_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output27 (.I(net27),
    .Z(data_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output28 (.I(net28),
    .Z(irq1));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output29 (.I(net29),
    .Z(irq2));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output30 (.I(net30),
    .Z(irq5));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output31 (.I(net31),
    .Z(pwm0));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output32 (.I(net32),
    .Z(pwm1));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output33 (.I(net33),
    .Z(pwm2));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output34 (.I(net34),
    .Z(tmr0_o));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output35 (.I(net35),
    .Z(tmr1_o));
endmodule

