magic
tech gf180mcuD
magscale 1 10
timestamp 1700749127
<< nwell >>
rect 1258 146176 148710 146694
rect 1258 145447 12776 145472
rect 1258 144633 148710 145447
rect 1258 144608 7581 144633
rect 1258 143879 3885 143904
rect 1258 143065 148710 143879
rect 1258 143040 2541 143065
rect 1258 142311 12440 142336
rect 1258 141497 148710 142311
rect 1258 141472 66760 141497
rect 1258 140743 18221 140768
rect 1258 139929 148710 140743
rect 1258 139904 2541 139929
rect 1258 139175 28413 139200
rect 1258 138361 148710 139175
rect 1258 138336 2541 138361
rect 1258 137607 21064 137632
rect 1258 136793 148710 137607
rect 1258 136768 29981 136793
rect 1258 136039 2541 136064
rect 1258 135225 148710 136039
rect 1258 135200 7870 135225
rect 1258 134471 4566 134496
rect 1258 133657 148710 134471
rect 1258 133632 16206 133657
rect 1258 132903 36029 132928
rect 1258 132089 148710 132903
rect 1258 132064 2998 132089
rect 1258 131335 7383 131360
rect 1258 130521 148710 131335
rect 1258 130496 7646 130521
rect 1258 129767 5182 129792
rect 1258 128953 148710 129767
rect 1258 128928 10334 128953
rect 1258 128199 28008 128224
rect 1258 127385 148710 128199
rect 1258 127360 2541 127385
rect 1258 126631 37192 126656
rect 1258 125817 148710 126631
rect 1258 125792 6461 125817
rect 1258 125063 2541 125088
rect 1258 124249 148710 125063
rect 1258 124224 10200 124249
rect 1258 123495 28904 123520
rect 1258 122681 148710 123495
rect 1258 122656 16718 122681
rect 1258 121927 3677 121952
rect 1258 121113 148710 121927
rect 1258 121088 4242 121113
rect 1258 120359 11286 120384
rect 1258 119545 148710 120359
rect 1258 119520 14991 119545
rect 1258 118791 7617 118816
rect 1258 117977 148710 118791
rect 1258 117952 16235 117977
rect 1258 117223 1999 117248
rect 1258 116409 148710 117223
rect 1258 116384 11062 116409
rect 1258 115655 27336 115680
rect 1258 114841 148710 115655
rect 1258 114816 7926 114841
rect 1258 114087 5406 114112
rect 1258 113273 148710 114087
rect 1258 113248 16046 113273
rect 1258 112519 11566 112544
rect 1258 111705 148710 112519
rect 1258 111680 40888 111705
rect 1258 110951 26173 110976
rect 1258 110137 148710 110951
rect 1258 110112 22141 110137
rect 1258 109383 44989 109408
rect 1258 108569 148710 109383
rect 1258 108544 9662 108569
rect 1258 107815 44541 107840
rect 1258 107001 148710 107815
rect 1258 106976 4398 107001
rect 1258 106247 30093 106272
rect 1258 105433 148710 106247
rect 1258 105408 40776 105433
rect 1258 104679 2541 104704
rect 1258 103865 148710 104679
rect 1258 103840 14301 103865
rect 1258 103111 3661 103136
rect 1258 102297 148710 103111
rect 1258 102272 2541 102297
rect 1258 101543 18557 101568
rect 1258 100729 148710 101543
rect 1258 100704 33005 100729
rect 1258 99975 6909 100000
rect 1258 99161 148710 99975
rect 1258 99136 17390 99161
rect 1258 98407 4221 98432
rect 1258 97593 148710 98407
rect 1258 97568 2541 97593
rect 1258 96839 28525 96864
rect 1258 96025 148710 96839
rect 1258 96000 31885 96025
rect 1258 95271 18148 95296
rect 1258 94457 148710 95271
rect 1258 94432 2541 94457
rect 1258 93703 10446 93728
rect 1258 92889 148710 93703
rect 1258 92864 8180 92889
rect 1258 92135 7823 92160
rect 1258 91321 148710 92135
rect 1258 91296 8495 91321
rect 1258 90567 34125 90592
rect 1258 89753 148710 90567
rect 1258 89728 2541 89753
rect 1258 88999 12303 89024
rect 1258 88185 148710 88999
rect 1258 88160 22141 88185
rect 1258 87431 22318 87456
rect 1258 86617 148710 87431
rect 1258 86592 16696 86617
rect 1258 85863 2541 85888
rect 1258 85049 148710 85863
rect 1258 85024 30765 85049
rect 1258 84295 11389 84320
rect 1258 83481 148710 84295
rect 1258 83456 37501 83481
rect 1258 82727 57421 82752
rect 1258 81913 148710 82727
rect 1258 81888 8378 81913
rect 1258 81159 2541 81184
rect 1258 80345 148710 81159
rect 1258 80320 30877 80345
rect 1258 79591 2541 79616
rect 1258 78777 148710 79591
rect 1258 78752 5802 78777
rect 1258 78023 7711 78048
rect 1258 77209 148710 78023
rect 1258 77184 7366 77209
rect 1258 76455 41853 76480
rect 1258 75641 148710 76455
rect 1258 75616 22477 75641
rect 1258 74887 2541 74912
rect 1258 74073 148710 74887
rect 1258 74048 15388 74073
rect 1258 73319 10572 73344
rect 1258 72505 148710 73319
rect 1258 72480 2653 72505
rect 1258 71751 22072 71776
rect 1258 70937 148710 71751
rect 1258 70912 41965 70937
rect 1258 70183 26014 70208
rect 1258 69369 148710 70183
rect 1258 69344 67061 69369
rect 1258 68615 2541 68640
rect 1258 67801 148710 68615
rect 1258 67776 2653 67801
rect 1258 67047 19677 67072
rect 1258 66233 148710 67047
rect 1258 66208 32152 66233
rect 1258 65479 43775 65504
rect 1258 64665 148710 65479
rect 1258 64640 17704 64665
rect 1258 63911 3213 63936
rect 1258 63097 148710 63911
rect 1258 63072 2541 63097
rect 1258 62343 6461 62368
rect 1258 61529 148710 62343
rect 1258 61504 18398 61529
rect 1258 60775 4893 60800
rect 1258 59961 148710 60775
rect 1258 59936 9149 59961
rect 1258 59207 12509 59232
rect 1258 58393 148710 59207
rect 1258 58368 8821 58393
rect 1258 57639 3390 57664
rect 1258 56825 148710 57639
rect 1258 56800 11804 56825
rect 1258 56071 10334 56096
rect 1258 55257 148710 56071
rect 1258 55232 29981 55257
rect 1258 54503 7275 54528
rect 1258 53689 148710 54503
rect 1258 53664 31852 53689
rect 1258 52935 51291 52960
rect 1258 52121 148710 52935
rect 1258 52096 40238 52121
rect 1258 51367 5910 51392
rect 1258 50553 148710 51367
rect 1258 50528 1990 50553
rect 1258 49799 33242 49824
rect 1258 48985 148710 49799
rect 1258 48960 31773 48985
rect 1258 48231 7590 48256
rect 1258 47417 148710 48231
rect 1258 47392 30930 47417
rect 1258 46663 10334 46688
rect 1258 45849 148710 46663
rect 1258 45824 42086 45849
rect 1258 45095 9718 45120
rect 1258 44281 148710 45095
rect 1258 44256 12574 44281
rect 1258 43527 82798 43552
rect 1258 42713 148710 43527
rect 1258 42688 45455 42713
rect 1258 41959 37382 41984
rect 1258 41145 148710 41959
rect 1258 41120 17278 41145
rect 1258 40391 27750 40416
rect 1258 39577 148710 40391
rect 1258 39552 8374 39577
rect 1258 38823 23718 38848
rect 1258 38009 148710 38823
rect 1258 37984 35478 38009
rect 1258 37255 2335 37280
rect 1258 36441 148710 37255
rect 1258 36416 5798 36441
rect 1258 35687 17901 35712
rect 1258 34873 148710 35687
rect 1258 34848 13638 34873
rect 1258 34119 4566 34144
rect 1258 33305 148710 34119
rect 1258 33280 49198 33305
rect 1258 32551 51887 32576
rect 1258 31737 148710 32551
rect 1258 31712 2550 31737
rect 1258 30983 1887 31008
rect 1258 30169 148710 30983
rect 1258 30144 9494 30169
rect 1258 29415 13526 29440
rect 1258 28601 148710 29415
rect 1258 28576 10278 28601
rect 1258 27847 52110 27872
rect 1258 27033 148710 27847
rect 1258 27008 11958 27033
rect 1258 26279 15878 26304
rect 1258 25465 148710 26279
rect 1258 25440 3670 25465
rect 1258 24711 7198 24736
rect 1258 23897 148710 24711
rect 1258 23872 6358 23897
rect 1258 23143 2998 23168
rect 1258 22329 148710 23143
rect 1258 22304 8108 22329
rect 1258 21575 3292 21600
rect 1258 20761 148710 21575
rect 1258 20736 6750 20761
rect 1258 20007 2998 20032
rect 1258 19193 148710 20007
rect 1258 19168 21590 19193
rect 1258 18439 6470 18464
rect 1258 17625 148710 18439
rect 1258 17600 4734 17625
rect 1258 16871 10460 16896
rect 1258 16057 148710 16871
rect 1258 16032 10173 16057
rect 1258 15303 8654 15328
rect 1258 14489 148710 15303
rect 1258 14464 10287 14489
rect 1258 13735 7198 13760
rect 1258 12921 148710 13735
rect 1258 12896 31455 12921
rect 1258 12167 10936 12192
rect 1258 11353 148710 12167
rect 1258 11328 13638 11353
rect 1258 10599 8654 10624
rect 1258 9785 148710 10599
rect 1258 9760 14991 9785
rect 1258 9031 10334 9056
rect 1258 8217 148710 9031
rect 1258 8192 22157 8217
rect 1258 7463 12518 7488
rect 1258 6649 148710 7463
rect 1258 6624 24684 6649
rect 1258 5895 15262 5920
rect 1258 5081 148710 5895
rect 1258 5056 23326 5081
rect 1258 4327 38738 4352
rect 1258 3488 148710 4327
<< pwell >>
rect 1258 145472 148710 146176
rect 1258 143904 148710 144608
rect 1258 142336 148710 143040
rect 1258 140768 148710 141472
rect 1258 139200 148710 139904
rect 1258 137632 148710 138336
rect 1258 136064 148710 136768
rect 1258 134496 148710 135200
rect 1258 132928 148710 133632
rect 1258 131360 148710 132064
rect 1258 129792 148710 130496
rect 1258 128224 148710 128928
rect 1258 126656 148710 127360
rect 1258 125088 148710 125792
rect 1258 123520 148710 124224
rect 1258 121952 148710 122656
rect 1258 120384 148710 121088
rect 1258 118816 148710 119520
rect 1258 117248 148710 117952
rect 1258 115680 148710 116384
rect 1258 114112 148710 114816
rect 1258 112544 148710 113248
rect 1258 110976 148710 111680
rect 1258 109408 148710 110112
rect 1258 107840 148710 108544
rect 1258 106272 148710 106976
rect 1258 104704 148710 105408
rect 1258 103136 148710 103840
rect 1258 101568 148710 102272
rect 1258 100000 148710 100704
rect 1258 98432 148710 99136
rect 1258 96864 148710 97568
rect 1258 95296 148710 96000
rect 1258 93728 148710 94432
rect 1258 92160 148710 92864
rect 1258 90592 148710 91296
rect 1258 89024 148710 89728
rect 1258 87456 148710 88160
rect 1258 85888 148710 86592
rect 1258 84320 148710 85024
rect 1258 82752 148710 83456
rect 1258 81184 148710 81888
rect 1258 79616 148710 80320
rect 1258 78048 148710 78752
rect 1258 76480 148710 77184
rect 1258 74912 148710 75616
rect 1258 73344 148710 74048
rect 1258 71776 148710 72480
rect 1258 70208 148710 70912
rect 1258 68640 148710 69344
rect 1258 67072 148710 67776
rect 1258 65504 148710 66208
rect 1258 63936 148710 64640
rect 1258 62368 148710 63072
rect 1258 60800 148710 61504
rect 1258 59232 148710 59936
rect 1258 57664 148710 58368
rect 1258 56096 148710 56800
rect 1258 54528 148710 55232
rect 1258 52960 148710 53664
rect 1258 51392 148710 52096
rect 1258 49824 148710 50528
rect 1258 48256 148710 48960
rect 1258 46688 148710 47392
rect 1258 45120 148710 45824
rect 1258 43552 148710 44256
rect 1258 41984 148710 42688
rect 1258 40416 148710 41120
rect 1258 38848 148710 39552
rect 1258 37280 148710 37984
rect 1258 35712 148710 36416
rect 1258 34144 148710 34848
rect 1258 32576 148710 33280
rect 1258 31008 148710 31712
rect 1258 29440 148710 30144
rect 1258 27872 148710 28576
rect 1258 26304 148710 27008
rect 1258 24736 148710 25440
rect 1258 23168 148710 23872
rect 1258 21600 148710 22304
rect 1258 20032 148710 20736
rect 1258 18464 148710 19168
rect 1258 16896 148710 17600
rect 1258 15328 148710 16032
rect 1258 13760 148710 14464
rect 1258 12192 148710 12896
rect 1258 10624 148710 11328
rect 1258 9056 148710 9760
rect 1258 7488 148710 8192
rect 1258 5920 148710 6624
rect 1258 4352 148710 5056
rect 1258 3050 148710 3488
<< obsm1 >>
rect 1344 3076 148624 146914
<< metal2 >>
rect 2688 149200 2800 150000
rect 7840 149200 7952 150000
rect 12992 149200 13104 150000
rect 18144 149200 18256 150000
rect 23296 149200 23408 150000
rect 28448 149200 28560 150000
rect 33600 149200 33712 150000
rect 38752 149200 38864 150000
rect 43904 149200 44016 150000
rect 49056 149200 49168 150000
rect 54208 149200 54320 150000
rect 59360 149200 59472 150000
rect 64512 149200 64624 150000
rect 69664 149200 69776 150000
rect 74816 149200 74928 150000
rect 79968 149200 80080 150000
rect 85120 149200 85232 150000
rect 90272 149200 90384 150000
rect 95424 149200 95536 150000
rect 100576 149200 100688 150000
rect 105728 149200 105840 150000
rect 110880 149200 110992 150000
rect 116032 149200 116144 150000
rect 121184 149200 121296 150000
rect 126336 149200 126448 150000
rect 131488 149200 131600 150000
rect 136640 149200 136752 150000
rect 141792 149200 141904 150000
rect 146944 149200 147056 150000
<< obsm2 >>
rect 1372 149140 2628 149200
rect 2860 149140 7780 149200
rect 8012 149140 12932 149200
rect 13164 149140 18084 149200
rect 18316 149140 23236 149200
rect 23468 149140 28388 149200
rect 28620 149140 33540 149200
rect 33772 149140 38692 149200
rect 38924 149140 43844 149200
rect 44076 149140 48996 149200
rect 49228 149140 54148 149200
rect 54380 149140 59300 149200
rect 59532 149140 64452 149200
rect 64684 149140 69604 149200
rect 69836 149140 74756 149200
rect 74988 149140 79908 149200
rect 80140 149140 85060 149200
rect 85292 149140 90212 149200
rect 90444 149140 95364 149200
rect 95596 149140 100516 149200
rect 100748 149140 105668 149200
rect 105900 149140 110820 149200
rect 111052 149140 115972 149200
rect 116204 149140 121124 149200
rect 121356 149140 126276 149200
rect 126508 149140 131428 149200
rect 131660 149140 136580 149200
rect 136812 149140 141732 149200
rect 141964 149140 146884 149200
rect 147116 149140 148260 149200
rect 1372 1474 148260 149140
<< obsm3 >>
rect 1362 1484 148270 146636
<< metal4 >>
rect 4448 3076 4768 146668
rect 19808 3076 20128 146668
rect 35168 3076 35488 146668
rect 50528 3076 50848 146668
rect 65888 3076 66208 146668
rect 81248 3076 81568 146668
rect 96608 3076 96928 146668
rect 111968 3076 112288 146668
rect 127328 3076 127648 146668
rect 142688 3076 143008 146668
<< obsm4 >>
rect 4284 3016 4388 146254
rect 4828 3016 19748 146254
rect 20188 3016 35108 146254
rect 35548 3016 50468 146254
rect 50908 3016 65828 146254
rect 66268 3016 81188 146254
rect 81628 3016 96548 146254
rect 96988 3016 111908 146254
rect 112348 3016 127268 146254
rect 127708 3016 141988 146254
rect 4284 1586 141988 3016
<< labels >>
rlabel metal2 s 2688 149200 2800 150000 6 DAC_clk
port 1 nsew signal output
rlabel metal2 s 12992 149200 13104 150000 6 DAC_dat_1
port 2 nsew signal output
rlabel metal2 s 18144 149200 18256 150000 6 DAC_dat_2
port 3 nsew signal output
rlabel metal2 s 7840 149200 7952 150000 6 DAC_le
port 4 nsew signal output
rlabel metal2 s 23296 149200 23408 150000 6 addr[0]
port 5 nsew signal input
rlabel metal2 s 28448 149200 28560 150000 6 addr[1]
port 6 nsew signal input
rlabel metal2 s 33600 149200 33712 150000 6 addr[2]
port 7 nsew signal input
rlabel metal2 s 38752 149200 38864 150000 6 addr[3]
port 8 nsew signal input
rlabel metal2 s 43904 149200 44016 150000 6 addr[4]
port 9 nsew signal input
rlabel metal2 s 131488 149200 131600 150000 6 bus_cyc
port 10 nsew signal input
rlabel metal2 s 49056 149200 49168 150000 6 bus_in[0]
port 11 nsew signal input
rlabel metal2 s 54208 149200 54320 150000 6 bus_in[1]
port 12 nsew signal input
rlabel metal2 s 59360 149200 59472 150000 6 bus_in[2]
port 13 nsew signal input
rlabel metal2 s 64512 149200 64624 150000 6 bus_in[3]
port 14 nsew signal input
rlabel metal2 s 69664 149200 69776 150000 6 bus_in[4]
port 15 nsew signal input
rlabel metal2 s 74816 149200 74928 150000 6 bus_in[5]
port 16 nsew signal input
rlabel metal2 s 79968 149200 80080 150000 6 bus_in[6]
port 17 nsew signal input
rlabel metal2 s 85120 149200 85232 150000 6 bus_in[7]
port 18 nsew signal input
rlabel metal2 s 90272 149200 90384 150000 6 bus_out[0]
port 19 nsew signal output
rlabel metal2 s 95424 149200 95536 150000 6 bus_out[1]
port 20 nsew signal output
rlabel metal2 s 100576 149200 100688 150000 6 bus_out[2]
port 21 nsew signal output
rlabel metal2 s 105728 149200 105840 150000 6 bus_out[3]
port 22 nsew signal output
rlabel metal2 s 110880 149200 110992 150000 6 bus_out[4]
port 23 nsew signal output
rlabel metal2 s 116032 149200 116144 150000 6 bus_out[5]
port 24 nsew signal output
rlabel metal2 s 121184 149200 121296 150000 6 bus_out[6]
port 25 nsew signal output
rlabel metal2 s 126336 149200 126448 150000 6 bus_out[7]
port 26 nsew signal output
rlabel metal2 s 136640 149200 136752 150000 6 bus_we
port 27 nsew signal input
rlabel metal2 s 141792 149200 141904 150000 6 clk
port 28 nsew signal input
rlabel metal2 s 146944 149200 147056 150000 6 rst
port 29 nsew signal input
rlabel metal4 s 4448 3076 4768 146668 6 vdd
port 30 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 146668 6 vdd
port 30 nsew power bidirectional
rlabel metal4 s 65888 3076 66208 146668 6 vdd
port 30 nsew power bidirectional
rlabel metal4 s 96608 3076 96928 146668 6 vdd
port 30 nsew power bidirectional
rlabel metal4 s 127328 3076 127648 146668 6 vdd
port 30 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 146668 6 vss
port 31 nsew ground bidirectional
rlabel metal4 s 50528 3076 50848 146668 6 vss
port 31 nsew ground bidirectional
rlabel metal4 s 81248 3076 81568 146668 6 vss
port 31 nsew ground bidirectional
rlabel metal4 s 111968 3076 112288 146668 6 vss
port 31 nsew ground bidirectional
rlabel metal4 s 142688 3076 143008 146668 6 vss
port 31 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 150000 150000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 17199140
string GDS_FILE /run/media/tholin/d9eb5833-69bc-462f-98fb-b7c5c019399b/AS2650/openlane/SID/runs/23_11_23_14_59/results/signoff/sid_top.magic.gds
string GDS_START 551084
<< end >>

