// This is the unpowered netlist.
module wrapped_as2650 (wb_clk_i,
    io_in,
    io_oeb,
    io_out);
 input wb_clk_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire _4300_;
 wire _4301_;
 wire _4302_;
 wire _4303_;
 wire _4304_;
 wire _4305_;
 wire _4306_;
 wire _4307_;
 wire _4308_;
 wire _4309_;
 wire _4310_;
 wire _4311_;
 wire _4312_;
 wire _4313_;
 wire _4314_;
 wire _4315_;
 wire _4316_;
 wire _4317_;
 wire _4318_;
 wire _4319_;
 wire _4320_;
 wire _4321_;
 wire _4322_;
 wire _4323_;
 wire _4324_;
 wire _4325_;
 wire _4326_;
 wire _4327_;
 wire _4328_;
 wire _4329_;
 wire _4330_;
 wire _4331_;
 wire _4332_;
 wire _4333_;
 wire _4334_;
 wire _4335_;
 wire _4336_;
 wire _4337_;
 wire _4338_;
 wire _4339_;
 wire _4340_;
 wire _4341_;
 wire _4342_;
 wire _4343_;
 wire _4344_;
 wire _4345_;
 wire _4346_;
 wire _4347_;
 wire _4348_;
 wire _4349_;
 wire _4350_;
 wire _4351_;
 wire _4352_;
 wire _4353_;
 wire _4354_;
 wire _4355_;
 wire _4356_;
 wire _4357_;
 wire _4358_;
 wire _4359_;
 wire _4360_;
 wire _4361_;
 wire _4362_;
 wire _4363_;
 wire _4364_;
 wire _4365_;
 wire _4366_;
 wire _4367_;
 wire _4368_;
 wire _4369_;
 wire _4370_;
 wire _4371_;
 wire _4372_;
 wire _4373_;
 wire _4374_;
 wire _4375_;
 wire _4376_;
 wire _4377_;
 wire _4378_;
 wire _4379_;
 wire _4380_;
 wire _4381_;
 wire _4382_;
 wire _4383_;
 wire _4384_;
 wire _4385_;
 wire _4386_;
 wire _4387_;
 wire _4388_;
 wire _4389_;
 wire _4390_;
 wire _4391_;
 wire _4392_;
 wire _4393_;
 wire _4394_;
 wire _4395_;
 wire _4396_;
 wire _4397_;
 wire _4398_;
 wire _4399_;
 wire _4400_;
 wire _4401_;
 wire _4402_;
 wire _4403_;
 wire _4404_;
 wire _4405_;
 wire _4406_;
 wire _4407_;
 wire _4408_;
 wire _4409_;
 wire _4410_;
 wire _4411_;
 wire _4412_;
 wire _4413_;
 wire _4414_;
 wire _4415_;
 wire _4416_;
 wire _4417_;
 wire _4418_;
 wire _4419_;
 wire _4420_;
 wire _4421_;
 wire _4422_;
 wire _4423_;
 wire _4424_;
 wire _4425_;
 wire _4426_;
 wire _4427_;
 wire _4428_;
 wire _4429_;
 wire _4430_;
 wire _4431_;
 wire _4432_;
 wire _4433_;
 wire _4434_;
 wire _4435_;
 wire _4436_;
 wire _4437_;
 wire _4438_;
 wire _4439_;
 wire _4440_;
 wire _4441_;
 wire _4442_;
 wire _4443_;
 wire _4444_;
 wire _4445_;
 wire _4446_;
 wire _4447_;
 wire _4448_;
 wire _4449_;
 wire _4450_;
 wire _4451_;
 wire _4452_;
 wire _4453_;
 wire _4454_;
 wire _4455_;
 wire _4456_;
 wire _4457_;
 wire _4458_;
 wire _4459_;
 wire _4460_;
 wire _4461_;
 wire _4462_;
 wire _4463_;
 wire _4464_;
 wire _4465_;
 wire _4466_;
 wire _4467_;
 wire _4468_;
 wire _4469_;
 wire _4470_;
 wire _4471_;
 wire _4472_;
 wire _4473_;
 wire _4474_;
 wire _4475_;
 wire _4476_;
 wire _4477_;
 wire _4478_;
 wire _4479_;
 wire _4480_;
 wire _4481_;
 wire _4482_;
 wire _4483_;
 wire _4484_;
 wire _4485_;
 wire _4486_;
 wire _4487_;
 wire _4488_;
 wire _4489_;
 wire _4490_;
 wire _4491_;
 wire _4492_;
 wire _4493_;
 wire _4494_;
 wire _4495_;
 wire _4496_;
 wire _4497_;
 wire _4498_;
 wire _4499_;
 wire _4500_;
 wire _4501_;
 wire _4502_;
 wire _4503_;
 wire _4504_;
 wire _4505_;
 wire _4506_;
 wire _4507_;
 wire _4508_;
 wire _4509_;
 wire _4510_;
 wire _4511_;
 wire _4512_;
 wire _4513_;
 wire _4514_;
 wire _4515_;
 wire _4516_;
 wire _4517_;
 wire _4518_;
 wire _4519_;
 wire _4520_;
 wire _4521_;
 wire _4522_;
 wire _4523_;
 wire _4524_;
 wire \as2650.addr_buff[0] ;
 wire \as2650.addr_buff[1] ;
 wire \as2650.addr_buff[2] ;
 wire \as2650.addr_buff[3] ;
 wire \as2650.addr_buff[4] ;
 wire \as2650.addr_buff[5] ;
 wire \as2650.addr_buff[6] ;
 wire \as2650.addr_buff[7] ;
 wire \as2650.alu_op[0] ;
 wire \as2650.alu_op[1] ;
 wire \as2650.alu_op[2] ;
 wire \as2650.carry ;
 wire \as2650.cycle[0] ;
 wire \as2650.cycle[1] ;
 wire \as2650.cycle[2] ;
 wire \as2650.cycle[3] ;
 wire \as2650.cycle[4] ;
 wire \as2650.cycle[5] ;
 wire \as2650.cycle[6] ;
 wire \as2650.cycle[7] ;
 wire \as2650.halted ;
 wire \as2650.holding_reg[0] ;
 wire \as2650.holding_reg[1] ;
 wire \as2650.holding_reg[2] ;
 wire \as2650.holding_reg[3] ;
 wire \as2650.holding_reg[4] ;
 wire \as2650.holding_reg[5] ;
 wire \as2650.holding_reg[6] ;
 wire \as2650.holding_reg[7] ;
 wire \as2650.idx_ctrl[0] ;
 wire \as2650.idx_ctrl[1] ;
 wire \as2650.ins_reg[0] ;
 wire \as2650.ins_reg[1] ;
 wire \as2650.ins_reg[2] ;
 wire \as2650.ins_reg[3] ;
 wire \as2650.ins_reg[4] ;
 wire \as2650.overflow ;
 wire \as2650.pc[0] ;
 wire \as2650.pc[10] ;
 wire \as2650.pc[11] ;
 wire \as2650.pc[12] ;
 wire \as2650.pc[13] ;
 wire \as2650.pc[14] ;
 wire \as2650.pc[1] ;
 wire \as2650.pc[2] ;
 wire \as2650.pc[3] ;
 wire \as2650.pc[4] ;
 wire \as2650.pc[5] ;
 wire \as2650.pc[6] ;
 wire \as2650.pc[7] ;
 wire \as2650.pc[8] ;
 wire \as2650.pc[9] ;
 wire \as2650.psl[1] ;
 wire \as2650.psl[3] ;
 wire \as2650.psl[4] ;
 wire \as2650.psl[5] ;
 wire \as2650.psl[6] ;
 wire \as2650.psl[7] ;
 wire \as2650.psu[0] ;
 wire \as2650.psu[1] ;
 wire \as2650.psu[2] ;
 wire \as2650.psu[3] ;
 wire \as2650.psu[4] ;
 wire \as2650.psu[5] ;
 wire \as2650.psu[7] ;
 wire \as2650.r0[0] ;
 wire \as2650.r0[1] ;
 wire \as2650.r0[2] ;
 wire \as2650.r0[3] ;
 wire \as2650.r0[4] ;
 wire \as2650.r0[5] ;
 wire \as2650.r0[6] ;
 wire \as2650.r0[7] ;
 wire \as2650.r123[0][0] ;
 wire \as2650.r123[0][1] ;
 wire \as2650.r123[0][2] ;
 wire \as2650.r123[0][3] ;
 wire \as2650.r123[0][4] ;
 wire \as2650.r123[0][5] ;
 wire \as2650.r123[0][6] ;
 wire \as2650.r123[0][7] ;
 wire \as2650.r123[1][0] ;
 wire \as2650.r123[1][1] ;
 wire \as2650.r123[1][2] ;
 wire \as2650.r123[1][3] ;
 wire \as2650.r123[1][4] ;
 wire \as2650.r123[1][5] ;
 wire \as2650.r123[1][6] ;
 wire \as2650.r123[1][7] ;
 wire \as2650.r123[2][0] ;
 wire \as2650.r123[2][1] ;
 wire \as2650.r123[2][2] ;
 wire \as2650.r123[2][3] ;
 wire \as2650.r123[2][4] ;
 wire \as2650.r123[2][5] ;
 wire \as2650.r123[2][6] ;
 wire \as2650.r123[2][7] ;
 wire \as2650.r123[3][0] ;
 wire \as2650.r123[3][1] ;
 wire \as2650.r123[3][2] ;
 wire \as2650.r123[3][3] ;
 wire \as2650.r123[3][4] ;
 wire \as2650.r123[3][5] ;
 wire \as2650.r123[3][6] ;
 wire \as2650.r123[3][7] ;
 wire \as2650.r123_2[0][0] ;
 wire \as2650.r123_2[0][1] ;
 wire \as2650.r123_2[0][2] ;
 wire \as2650.r123_2[0][3] ;
 wire \as2650.r123_2[0][4] ;
 wire \as2650.r123_2[0][5] ;
 wire \as2650.r123_2[0][6] ;
 wire \as2650.r123_2[0][7] ;
 wire \as2650.r123_2[1][0] ;
 wire \as2650.r123_2[1][1] ;
 wire \as2650.r123_2[1][2] ;
 wire \as2650.r123_2[1][3] ;
 wire \as2650.r123_2[1][4] ;
 wire \as2650.r123_2[1][5] ;
 wire \as2650.r123_2[1][6] ;
 wire \as2650.r123_2[1][7] ;
 wire \as2650.r123_2[2][0] ;
 wire \as2650.r123_2[2][1] ;
 wire \as2650.r123_2[2][2] ;
 wire \as2650.r123_2[2][3] ;
 wire \as2650.r123_2[2][4] ;
 wire \as2650.r123_2[2][5] ;
 wire \as2650.r123_2[2][6] ;
 wire \as2650.r123_2[2][7] ;
 wire \as2650.r123_2[3][0] ;
 wire \as2650.r123_2[3][1] ;
 wire \as2650.r123_2[3][2] ;
 wire \as2650.r123_2[3][3] ;
 wire \as2650.r123_2[3][4] ;
 wire \as2650.r123_2[3][5] ;
 wire \as2650.r123_2[3][6] ;
 wire \as2650.r123_2[3][7] ;
 wire \as2650.stack[0][0] ;
 wire \as2650.stack[0][10] ;
 wire \as2650.stack[0][11] ;
 wire \as2650.stack[0][12] ;
 wire \as2650.stack[0][13] ;
 wire \as2650.stack[0][14] ;
 wire \as2650.stack[0][1] ;
 wire \as2650.stack[0][2] ;
 wire \as2650.stack[0][3] ;
 wire \as2650.stack[0][4] ;
 wire \as2650.stack[0][5] ;
 wire \as2650.stack[0][6] ;
 wire \as2650.stack[0][7] ;
 wire \as2650.stack[0][8] ;
 wire \as2650.stack[0][9] ;
 wire \as2650.stack[1][0] ;
 wire \as2650.stack[1][10] ;
 wire \as2650.stack[1][11] ;
 wire \as2650.stack[1][12] ;
 wire \as2650.stack[1][13] ;
 wire \as2650.stack[1][14] ;
 wire \as2650.stack[1][1] ;
 wire \as2650.stack[1][2] ;
 wire \as2650.stack[1][3] ;
 wire \as2650.stack[1][4] ;
 wire \as2650.stack[1][5] ;
 wire \as2650.stack[1][6] ;
 wire \as2650.stack[1][7] ;
 wire \as2650.stack[1][8] ;
 wire \as2650.stack[1][9] ;
 wire \as2650.stack[2][0] ;
 wire \as2650.stack[2][10] ;
 wire \as2650.stack[2][11] ;
 wire \as2650.stack[2][12] ;
 wire \as2650.stack[2][13] ;
 wire \as2650.stack[2][14] ;
 wire \as2650.stack[2][1] ;
 wire \as2650.stack[2][2] ;
 wire \as2650.stack[2][3] ;
 wire \as2650.stack[2][4] ;
 wire \as2650.stack[2][5] ;
 wire \as2650.stack[2][6] ;
 wire \as2650.stack[2][7] ;
 wire \as2650.stack[2][8] ;
 wire \as2650.stack[2][9] ;
 wire \as2650.stack[3][0] ;
 wire \as2650.stack[3][10] ;
 wire \as2650.stack[3][11] ;
 wire \as2650.stack[3][12] ;
 wire \as2650.stack[3][13] ;
 wire \as2650.stack[3][14] ;
 wire \as2650.stack[3][1] ;
 wire \as2650.stack[3][2] ;
 wire \as2650.stack[3][3] ;
 wire \as2650.stack[3][4] ;
 wire \as2650.stack[3][5] ;
 wire \as2650.stack[3][6] ;
 wire \as2650.stack[3][7] ;
 wire \as2650.stack[3][8] ;
 wire \as2650.stack[3][9] ;
 wire \as2650.stack[4][0] ;
 wire \as2650.stack[4][10] ;
 wire \as2650.stack[4][11] ;
 wire \as2650.stack[4][12] ;
 wire \as2650.stack[4][13] ;
 wire \as2650.stack[4][14] ;
 wire \as2650.stack[4][1] ;
 wire \as2650.stack[4][2] ;
 wire \as2650.stack[4][3] ;
 wire \as2650.stack[4][4] ;
 wire \as2650.stack[4][5] ;
 wire \as2650.stack[4][6] ;
 wire \as2650.stack[4][7] ;
 wire \as2650.stack[4][8] ;
 wire \as2650.stack[4][9] ;
 wire \as2650.stack[5][0] ;
 wire \as2650.stack[5][10] ;
 wire \as2650.stack[5][11] ;
 wire \as2650.stack[5][12] ;
 wire \as2650.stack[5][13] ;
 wire \as2650.stack[5][14] ;
 wire \as2650.stack[5][1] ;
 wire \as2650.stack[5][2] ;
 wire \as2650.stack[5][3] ;
 wire \as2650.stack[5][4] ;
 wire \as2650.stack[5][5] ;
 wire \as2650.stack[5][6] ;
 wire \as2650.stack[5][7] ;
 wire \as2650.stack[5][8] ;
 wire \as2650.stack[5][9] ;
 wire \as2650.stack[6][0] ;
 wire \as2650.stack[6][10] ;
 wire \as2650.stack[6][11] ;
 wire \as2650.stack[6][12] ;
 wire \as2650.stack[6][13] ;
 wire \as2650.stack[6][14] ;
 wire \as2650.stack[6][1] ;
 wire \as2650.stack[6][2] ;
 wire \as2650.stack[6][3] ;
 wire \as2650.stack[6][4] ;
 wire \as2650.stack[6][5] ;
 wire \as2650.stack[6][6] ;
 wire \as2650.stack[6][7] ;
 wire \as2650.stack[6][8] ;
 wire \as2650.stack[6][9] ;
 wire \as2650.stack[7][0] ;
 wire \as2650.stack[7][10] ;
 wire \as2650.stack[7][11] ;
 wire \as2650.stack[7][12] ;
 wire \as2650.stack[7][13] ;
 wire \as2650.stack[7][14] ;
 wire \as2650.stack[7][1] ;
 wire \as2650.stack[7][2] ;
 wire \as2650.stack[7][3] ;
 wire \as2650.stack[7][4] ;
 wire \as2650.stack[7][5] ;
 wire \as2650.stack[7][6] ;
 wire \as2650.stack[7][7] ;
 wire \as2650.stack[7][8] ;
 wire \as2650.stack[7][9] ;
 wire net86;
 wire net91;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net87;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net88;
 wire net72;
 wire net73;
 wire net74;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire clknet_leaf_0_wb_clk_i;
 wire net89;
 wire net90;
 wire net75;
 wire net80;
 wire net76;
 wire net77;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net78;
 wire net79;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_57_wb_clk_i;
 wire clknet_leaf_58_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_60_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_62_wb_clk_i;
 wire clknet_leaf_63_wb_clk_i;
 wire clknet_leaf_65_wb_clk_i;
 wire clknet_leaf_66_wb_clk_i;
 wire clknet_leaf_67_wb_clk_i;
 wire clknet_leaf_68_wb_clk_i;
 wire clknet_leaf_69_wb_clk_i;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0__leaf_wb_clk_i;
 wire clknet_3_1__leaf_wb_clk_i;
 wire clknet_3_2__leaf_wb_clk_i;
 wire clknet_3_3__leaf_wb_clk_i;
 wire clknet_3_4__leaf_wb_clk_i;
 wire clknet_3_5__leaf_wb_clk_i;
 wire clknet_3_6__leaf_wb_clk_i;
 wire clknet_3_7__leaf_wb_clk_i;
 wire clknet_opt_1_0_wb_clk_i;
 wire clknet_opt_2_0_wb_clk_i;
 wire clknet_opt_3_0_wb_clk_i;
 wire clknet_opt_4_0_wb_clk_i;
 wire clknet_opt_5_0_wb_clk_i;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4525_ (.I(net50),
    .ZN(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4526_ (.I(\as2650.r123[0][0] ),
    .ZN(_4107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4527_ (.I(\as2650.psl[4] ),
    .Z(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4528_ (.I(_4108_),
    .Z(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4529_ (.I(_4109_),
    .Z(_4110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4530_ (.I(_4110_),
    .Z(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4531_ (.I(_4111_),
    .Z(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4532_ (.I(_4112_),
    .Z(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4533_ (.I(\as2650.halted ),
    .Z(_4114_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4534_ (.I(_4114_),
    .ZN(_4115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4535_ (.I(net5),
    .ZN(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4536_ (.A1(_4115_),
    .A2(_4116_),
    .ZN(_4117_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4537_ (.A1(_4113_),
    .A2(_4117_),
    .ZN(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4538_ (.I(\as2650.cycle[0] ),
    .Z(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4539_ (.I(\as2650.cycle[2] ),
    .Z(_4120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4540_ (.I(\as2650.cycle[5] ),
    .Z(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _4541_ (.A1(\as2650.cycle[7] ),
    .A2(\as2650.cycle[6] ),
    .A3(_4121_),
    .A4(\as2650.cycle[4] ),
    .Z(_4122_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4542_ (.A1(\as2650.cycle[3] ),
    .A2(_4120_),
    .A3(_4122_),
    .ZN(_4123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4543_ (.A1(\as2650.cycle[1] ),
    .A2(_4123_),
    .ZN(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4544_ (.A1(_4119_),
    .A2(_4124_),
    .ZN(_4125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4545_ (.I(_4125_),
    .Z(_4126_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4546_ (.A1(_4118_),
    .A2(_4126_),
    .Z(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4547_ (.I(\as2650.ins_reg[3] ),
    .Z(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4548_ (.A1(\as2650.ins_reg[2] ),
    .A2(_4128_),
    .ZN(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4549_ (.I(_4129_),
    .Z(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4550_ (.I(_4130_),
    .Z(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4551_ (.I(_4131_),
    .Z(_4132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4552_ (.I(_4132_),
    .Z(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4553_ (.I(\as2650.alu_op[0] ),
    .ZN(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4554_ (.I(_4134_),
    .Z(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4555_ (.I(\as2650.ins_reg[4] ),
    .Z(_4136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4556_ (.I(_4136_),
    .Z(_4137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4557_ (.A1(_4135_),
    .A2(_4137_),
    .ZN(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4558_ (.I(\as2650.alu_op[1] ),
    .Z(_4139_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4559_ (.I(_4139_),
    .ZN(_4140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4560_ (.I(_4140_),
    .Z(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4561_ (.I(\as2650.alu_op[2] ),
    .Z(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4562_ (.I(_4142_),
    .Z(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4563_ (.A1(_4141_),
    .A2(_4143_),
    .ZN(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4564_ (.A1(_4138_),
    .A2(_4144_),
    .ZN(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4565_ (.I(\as2650.ins_reg[0] ),
    .Z(_4146_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4566_ (.I(_4146_),
    .ZN(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4567_ (.I(_4147_),
    .Z(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4568_ (.I(\as2650.ins_reg[1] ),
    .Z(_4149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4569_ (.I(_4149_),
    .Z(_4150_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4570_ (.A1(_4148_),
    .A2(_4150_),
    .ZN(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4571_ (.A1(_4133_),
    .A2(_4145_),
    .A3(_4151_),
    .ZN(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4572_ (.I(\as2650.alu_op[0] ),
    .Z(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4573_ (.I(_4153_),
    .Z(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4574_ (.I(_4139_),
    .Z(_4155_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4575_ (.A1(_4155_),
    .A2(_4142_),
    .ZN(_4156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4576_ (.A1(_4137_),
    .A2(_4156_),
    .ZN(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4577_ (.A1(_4154_),
    .A2(_4157_),
    .ZN(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4578_ (.A1(\as2650.ins_reg[2] ),
    .A2(\as2650.ins_reg[3] ),
    .Z(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4579_ (.I(_4159_),
    .Z(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4580_ (.I(_4160_),
    .Z(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4581_ (.I(_4161_),
    .Z(_4162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4582_ (.I(_4162_),
    .Z(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4583_ (.I(_4149_),
    .ZN(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4584_ (.A1(_4148_),
    .A2(_4164_),
    .ZN(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4585_ (.I(_4165_),
    .Z(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4586_ (.A1(_4163_),
    .A2(_4166_),
    .ZN(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4587_ (.A1(_4158_),
    .A2(_4167_),
    .ZN(_4168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4588_ (.A1(_4152_),
    .A2(_4168_),
    .ZN(_4169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4589_ (.I(_4169_),
    .Z(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4590_ (.I(_4150_),
    .Z(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4591_ (.A1(\as2650.halted ),
    .A2(net5),
    .ZN(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4592_ (.I(\as2650.ins_reg[0] ),
    .Z(_4173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4593_ (.A1(_4173_),
    .A2(\as2650.ins_reg[1] ),
    .ZN(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4594_ (.I(_4174_),
    .Z(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4595_ (.I(_4175_),
    .Z(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4596_ (.I(_4176_),
    .Z(_4177_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4597_ (.A1(_4113_),
    .A2(_4177_),
    .ZN(_4178_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4598_ (.A1(_4172_),
    .A2(_4178_),
    .Z(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4599_ (.I(_4179_),
    .Z(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4600_ (.I(_4137_),
    .Z(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4601_ (.I(_4181_),
    .Z(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4602_ (.A1(_4155_),
    .A2(_4182_),
    .ZN(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4603_ (.I(_4128_),
    .Z(_4184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4604_ (.I(_4184_),
    .Z(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4605_ (.I(_4126_),
    .Z(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4606_ (.A1(_4185_),
    .A2(_4186_),
    .ZN(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4607_ (.I(\as2650.cycle[3] ),
    .ZN(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4608_ (.I(\as2650.cycle[2] ),
    .ZN(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4609_ (.A1(\as2650.cycle[7] ),
    .A2(\as2650.cycle[6] ),
    .A3(\as2650.cycle[5] ),
    .A4(\as2650.cycle[4] ),
    .ZN(_4190_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4610_ (.A1(_4188_),
    .A2(_4189_),
    .A3(_4190_),
    .ZN(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4611_ (.I(\as2650.cycle[1] ),
    .Z(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4612_ (.I(\as2650.cycle[0] ),
    .Z(_4193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4613_ (.A1(_4192_),
    .A2(_4193_),
    .ZN(_4194_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4614_ (.A1(_4191_),
    .A2(_4194_),
    .ZN(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4615_ (.I(_4142_),
    .ZN(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4616_ (.I(\as2650.ins_reg[2] ),
    .Z(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4617_ (.I(_4136_),
    .Z(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4618_ (.A1(_4153_),
    .A2(_4198_),
    .ZN(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4619_ (.A1(_4197_),
    .A2(_4199_),
    .ZN(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4620_ (.A1(_4196_),
    .A2(_4200_),
    .ZN(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4621_ (.A1(_4184_),
    .A2(_4201_),
    .ZN(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4622_ (.A1(_4195_),
    .A2(_4202_),
    .ZN(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4623_ (.A1(_4183_),
    .A2(_4187_),
    .B(_4203_),
    .ZN(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4624_ (.A1(_4180_),
    .A2(_4204_),
    .Z(_4205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4625_ (.I(_4186_),
    .Z(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4626_ (.I(_4178_),
    .Z(_4207_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4627_ (.I(_4197_),
    .ZN(_4208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4628_ (.I(_4208_),
    .Z(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4629_ (.I(_4209_),
    .Z(_4210_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4630_ (.A1(_4139_),
    .A2(\as2650.alu_op[2] ),
    .A3(\as2650.ins_reg[4] ),
    .ZN(_4211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4631_ (.A1(\as2650.alu_op[0] ),
    .A2(_4211_),
    .ZN(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4632_ (.A1(_4210_),
    .A2(_4212_),
    .ZN(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4633_ (.A1(_4184_),
    .A2(_4117_),
    .A3(_4213_),
    .ZN(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4634_ (.A1(_4206_),
    .A2(_4207_),
    .A3(_4214_),
    .Z(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4635_ (.I(_4128_),
    .Z(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4636_ (.I(_4198_),
    .Z(_4217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4637_ (.A1(_4140_),
    .A2(_4142_),
    .ZN(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4638_ (.A1(_4209_),
    .A2(_4135_),
    .A3(_4217_),
    .A4(_4218_),
    .ZN(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4639_ (.A1(_4216_),
    .A2(_4219_),
    .ZN(_4220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4640_ (.I(_4125_),
    .Z(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4641_ (.I(_4221_),
    .Z(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4642_ (.A1(_4220_),
    .A2(_4222_),
    .A3(_4180_),
    .ZN(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4643_ (.I(_4221_),
    .Z(_4224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4644_ (.I(_4217_),
    .Z(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4645_ (.I(_4163_),
    .Z(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4646_ (.I(_4226_),
    .Z(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4647_ (.A1(_4155_),
    .A2(_4134_),
    .A3(_4143_),
    .ZN(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4648_ (.A1(_4225_),
    .A2(_4227_),
    .A3(_4228_),
    .ZN(_4229_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4649_ (.A1(_4224_),
    .A2(_4180_),
    .A3(_4229_),
    .ZN(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4650_ (.A1(_4223_),
    .A2(_4230_),
    .ZN(_4231_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4651_ (.I(_4137_),
    .ZN(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4652_ (.I(_4232_),
    .Z(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4653_ (.I(_4233_),
    .Z(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4654_ (.I(\as2650.cycle[7] ),
    .Z(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4655_ (.I(\as2650.cycle[1] ),
    .ZN(_4236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4656_ (.A1(_4236_),
    .A2(_4119_),
    .ZN(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4657_ (.I(\as2650.cycle[3] ),
    .Z(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4658_ (.A1(_4121_),
    .A2(\as2650.cycle[4] ),
    .A3(_4238_),
    .A4(_4120_),
    .ZN(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4659_ (.A1(\as2650.cycle[6] ),
    .A2(_4239_),
    .ZN(_4240_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4660_ (.A1(_4237_),
    .A2(_4240_),
    .ZN(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4661_ (.A1(_4235_),
    .A2(_4241_),
    .ZN(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4662_ (.I(\as2650.addr_buff[6] ),
    .Z(_4243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4663_ (.I(\as2650.addr_buff[5] ),
    .Z(_4244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4664_ (.A1(_4243_),
    .A2(_4244_),
    .ZN(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4665_ (.A1(\as2650.addr_buff[7] ),
    .A2(_4245_),
    .Z(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4666_ (.A1(_4242_),
    .A2(_4246_),
    .ZN(_4247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4667_ (.I(_4247_),
    .Z(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4668_ (.A1(_4234_),
    .A2(_4180_),
    .A3(_4248_),
    .ZN(_4249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4669_ (.I(_4181_),
    .Z(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4670_ (.I(_4250_),
    .Z(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4671_ (.A1(_4192_),
    .A2(_4119_),
    .ZN(_4252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4672_ (.A1(_4188_),
    .A2(_4120_),
    .ZN(_4253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4673_ (.A1(_4122_),
    .A2(_4253_),
    .ZN(_4254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4674_ (.A1(_4252_),
    .A2(_4254_),
    .ZN(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4675_ (.I(_4255_),
    .Z(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4676_ (.I(_4177_),
    .Z(_4257_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4677_ (.A1(\as2650.idx_ctrl[1] ),
    .A2(\as2650.idx_ctrl[0] ),
    .Z(_4258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4678_ (.I(_4258_),
    .Z(_4259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4679_ (.I(_4259_),
    .Z(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4680_ (.A1(\as2650.alu_op[1] ),
    .A2(\as2650.alu_op[2] ),
    .ZN(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4681_ (.A1(_4134_),
    .A2(_4261_),
    .ZN(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4682_ (.I(_4262_),
    .Z(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _4683_ (.A1(_4133_),
    .A2(_4257_),
    .A3(_4260_),
    .A4(_4263_),
    .Z(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4684_ (.A1(_4251_),
    .A2(_4256_),
    .A3(_4264_),
    .ZN(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4685_ (.A1(_4118_),
    .A2(_4265_),
    .ZN(_4266_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4686_ (.A1(_4237_),
    .A2(_4240_),
    .Z(_4267_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4687_ (.A1(_4235_),
    .A2(_4267_),
    .ZN(_4268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4688_ (.I(_4268_),
    .Z(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4689_ (.I(_4117_),
    .Z(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4690_ (.A1(_4250_),
    .A2(_4270_),
    .ZN(_4271_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4691_ (.I(_4271_),
    .ZN(_4272_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4692_ (.A1(\as2650.idx_ctrl[1] ),
    .A2(\as2650.idx_ctrl[0] ),
    .ZN(_4273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4693_ (.I(_4273_),
    .Z(_4274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4694_ (.I(_4274_),
    .Z(_4275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4695_ (.I(_4275_),
    .Z(_4276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4696_ (.I(_4276_),
    .Z(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4697_ (.I(_4277_),
    .Z(_4278_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4698_ (.A1(_4272_),
    .A2(_4278_),
    .ZN(_4279_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4699_ (.A1(_4207_),
    .A2(_4269_),
    .A3(_4279_),
    .ZN(_4280_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4700_ (.A1(_4249_),
    .A2(_4266_),
    .A3(_4280_),
    .ZN(_4281_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _4701_ (.A1(_4205_),
    .A2(_4215_),
    .A3(_4231_),
    .A4(_4281_),
    .ZN(_4282_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4702_ (.A1(_4171_),
    .A2(_4282_),
    .ZN(_4283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4703_ (.I(net5),
    .Z(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4704_ (.A1(_4127_),
    .A2(_4170_),
    .B(_4283_),
    .C(_4284_),
    .ZN(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4705_ (.I(_4285_),
    .Z(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4706_ (.I(_4286_),
    .Z(_4287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4707_ (.I(_4283_),
    .Z(_4288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4708_ (.I(_4266_),
    .Z(_4289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4709_ (.I(_4289_),
    .Z(_4290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4710_ (.A1(_4155_),
    .A2(_4196_),
    .ZN(_4291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4711_ (.I(_4291_),
    .Z(_4292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4712_ (.I(_4144_),
    .Z(_4293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4713_ (.I(_4156_),
    .Z(_4294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4714_ (.A1(_4154_),
    .A2(_4294_),
    .ZN(_4295_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4715_ (.A1(_4292_),
    .A2(_4293_),
    .A3(_4295_),
    .ZN(_4296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4716_ (.I(_4296_),
    .Z(_4297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4717_ (.I(_4297_),
    .Z(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4718_ (.I(\as2650.r0[0] ),
    .Z(_4299_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4719_ (.A1(_4146_),
    .A2(_4149_),
    .Z(_4300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4720_ (.I(_4110_),
    .Z(_4301_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4721_ (.I0(\as2650.r123[2][0] ),
    .I1(\as2650.r123_2[2][0] ),
    .S(_4301_),
    .Z(_4302_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4722_ (.A1(_4173_),
    .A2(\as2650.ins_reg[1] ),
    .Z(_4303_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4723_ (.I0(\as2650.r123[1][0] ),
    .I1(\as2650.r123[0][0] ),
    .I2(\as2650.r123_2[1][0] ),
    .I3(\as2650.r123_2[0][0] ),
    .S0(_4146_),
    .S1(_4301_),
    .Z(_4304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _4724_ (.A1(_4299_),
    .A2(_4175_),
    .B1(_4300_),
    .B2(_4302_),
    .C1(_4303_),
    .C2(_4304_),
    .ZN(_4305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4725_ (.I(_4305_),
    .Z(_4306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4726_ (.A1(\as2650.holding_reg[0] ),
    .A2(_4160_),
    .ZN(_4307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4727_ (.A1(_4160_),
    .A2(_4306_),
    .B(_4307_),
    .ZN(_4308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4728_ (.I(_4135_),
    .Z(_4309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4729_ (.I(_4309_),
    .Z(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4730_ (.I(_4310_),
    .Z(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4731_ (.A1(_4139_),
    .A2(_4196_),
    .ZN(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4732_ (.A1(_4311_),
    .A2(_4312_),
    .ZN(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4733_ (.A1(\as2650.psl[3] ),
    .A2(\as2650.carry ),
    .ZN(_4314_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4734_ (.I(_4314_),
    .ZN(_4315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4735_ (.I(_4299_),
    .Z(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4736_ (.I(_4316_),
    .Z(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4737_ (.A1(_4317_),
    .A2(_4258_),
    .ZN(_4318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4738_ (.I(_4159_),
    .Z(_4319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4739_ (.I(_4319_),
    .Z(_4320_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4740_ (.A1(_4259_),
    .A2(_4306_),
    .B(_4318_),
    .C(_4320_),
    .ZN(_4321_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4741_ (.I(\as2650.holding_reg[0] ),
    .ZN(_4322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4742_ (.I(_4129_),
    .Z(_4323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4743_ (.A1(_4322_),
    .A2(_4323_),
    .ZN(_4324_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4744_ (.A1(_4308_),
    .A2(_4321_),
    .A3(_4324_),
    .ZN(_4325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4745_ (.A1(_4317_),
    .A2(_4274_),
    .B(_4160_),
    .ZN(_4326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4746_ (.A1(_4274_),
    .A2(_4306_),
    .B(_4326_),
    .ZN(_4327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4747_ (.A1(_4322_),
    .A2(_4320_),
    .ZN(_4328_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4748_ (.A1(_4308_),
    .A2(_4327_),
    .A3(_4328_),
    .Z(_4329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4749_ (.A1(_4325_),
    .A2(_4329_),
    .ZN(_4330_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4750_ (.A1(_4315_),
    .A2(_4330_),
    .Z(_4331_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4751_ (.A1(_4309_),
    .A2(_4293_),
    .ZN(_4332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4752_ (.I(_4332_),
    .Z(_4333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4753_ (.I(_4333_),
    .Z(_4334_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4754_ (.I(\as2650.carry ),
    .ZN(_4335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4755_ (.A1(\as2650.psl[3] ),
    .A2(_4335_),
    .ZN(_4336_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4756_ (.A1(_4336_),
    .A2(_4330_),
    .Z(_4337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4757_ (.I(_4295_),
    .Z(_4338_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4758_ (.A1(_4308_),
    .A2(_4321_),
    .A3(_4324_),
    .Z(_4339_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4759_ (.A1(_4153_),
    .A2(_4291_),
    .ZN(_4340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4760_ (.I(_4340_),
    .Z(_4341_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4761_ (.A1(_4309_),
    .A2(_4292_),
    .ZN(_4342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4762_ (.A1(_4339_),
    .A2(_4341_),
    .B1(_4342_),
    .B2(_4329_),
    .ZN(_4343_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4763_ (.A1(_4338_),
    .A2(_4330_),
    .B(_4343_),
    .C(_4297_),
    .ZN(_4344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4764_ (.A1(_4334_),
    .A2(_4337_),
    .B(_4344_),
    .ZN(_4345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4765_ (.A1(_4313_),
    .A2(_4331_),
    .B(_4345_),
    .ZN(_4346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4766_ (.A1(_4298_),
    .A2(_4308_),
    .B(_4346_),
    .ZN(_4347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4767_ (.I(_4289_),
    .Z(_4348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4768_ (.I(_4280_),
    .Z(_4349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4769_ (.I(_4349_),
    .Z(_4350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4770_ (.I(_4249_),
    .Z(_4351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4771_ (.I(_4351_),
    .Z(_4352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4772_ (.I(_4317_),
    .Z(_4353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4773_ (.I(_4353_),
    .Z(_4354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4774_ (.I(_4230_),
    .Z(_4355_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4775_ (.A1(_4222_),
    .A2(_4207_),
    .A3(_4214_),
    .ZN(_4356_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4776_ (.I(\as2650.psl[3] ),
    .Z(_4357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4777_ (.I(\as2650.r0[7] ),
    .Z(_4358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4778_ (.I(_4358_),
    .Z(_4359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4779_ (.A1(_4359_),
    .A2(_4176_),
    .ZN(_4360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4780_ (.I(_4300_),
    .Z(_4361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4781_ (.I(_4361_),
    .Z(_4362_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4782_ (.I0(\as2650.r123[2][7] ),
    .I1(\as2650.r123_2[2][7] ),
    .S(_4112_),
    .Z(_4363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4783_ (.A1(_4362_),
    .A2(_4363_),
    .ZN(_4364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4784_ (.I(_4303_),
    .Z(_4365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4785_ (.I(_4173_),
    .Z(_4366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4786_ (.I(_4366_),
    .Z(_4367_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4787_ (.I0(\as2650.r123[1][7] ),
    .I1(\as2650.r123[0][7] ),
    .I2(\as2650.r123_2[1][7] ),
    .I3(\as2650.r123_2[0][7] ),
    .S0(_4367_),
    .S1(_4112_),
    .Z(_4368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4788_ (.A1(_4365_),
    .A2(_4368_),
    .ZN(_4369_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4789_ (.A1(_4360_),
    .A2(_4364_),
    .A3(_4369_),
    .ZN(_4370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4790_ (.A1(_4357_),
    .A2(_4370_),
    .B(_4336_),
    .ZN(_4371_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4791_ (.I(_4166_),
    .Z(_4372_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4792_ (.A1(_4220_),
    .A2(_4372_),
    .A3(_4127_),
    .ZN(_4373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4793_ (.I(_4373_),
    .Z(_4374_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4794_ (.I(_4109_),
    .Z(_4375_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4795_ (.I0(\as2650.r123[1][1] ),
    .I1(\as2650.r123[0][1] ),
    .I2(\as2650.r123_2[1][1] ),
    .I3(\as2650.r123_2[0][1] ),
    .S0(_4173_),
    .S1(_4375_),
    .Z(_4376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4796_ (.A1(_4303_),
    .A2(_4376_),
    .ZN(_4377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4797_ (.I(_4377_),
    .Z(_4378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4798_ (.I(\as2650.r0[1] ),
    .Z(_4379_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4799_ (.I0(\as2650.r123[2][1] ),
    .I1(\as2650.r123_2[2][1] ),
    .S(_4375_),
    .Z(_4380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4800_ (.A1(_4379_),
    .A2(_4174_),
    .B1(_4300_),
    .B2(_4380_),
    .ZN(_4381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4801_ (.I(_4381_),
    .Z(_4382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4802_ (.A1(_4378_),
    .A2(_4382_),
    .ZN(_4383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4803_ (.I(_4383_),
    .Z(_4384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4804_ (.I(_4373_),
    .Z(_4385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4805_ (.I(net6),
    .Z(_4386_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4806_ (.I(_4386_),
    .Z(_4387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4807_ (.A1(_4236_),
    .A2(_4191_),
    .ZN(_4388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4808_ (.A1(_4193_),
    .A2(_4388_),
    .ZN(_4389_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4809_ (.I(_4128_),
    .ZN(_4390_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4810_ (.A1(_4208_),
    .A2(_4153_),
    .A3(_4198_),
    .ZN(_4391_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4811_ (.A1(_4143_),
    .A2(_4391_),
    .ZN(_4392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4812_ (.A1(_4390_),
    .A2(_4392_),
    .ZN(_4393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4813_ (.A1(_4389_),
    .A2(_4393_),
    .ZN(_4394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4814_ (.A1(_4179_),
    .A2(_4394_),
    .ZN(_4395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4815_ (.I(_4395_),
    .Z(_4396_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4816_ (.I(_4305_),
    .Z(_4397_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4817_ (.I(_4397_),
    .ZN(_4398_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4818_ (.A1(_4211_),
    .A2(_4398_),
    .Z(_4399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4819_ (.A1(_4399_),
    .A2(_4395_),
    .ZN(_4400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4820_ (.A1(_4387_),
    .A2(_4396_),
    .B(_4400_),
    .ZN(_4401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4821_ (.A1(_4385_),
    .A2(_4401_),
    .ZN(_4402_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4822_ (.I(_4111_),
    .ZN(_4403_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4823_ (.I(_4119_),
    .ZN(_4404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4824_ (.I(_4388_),
    .Z(_4405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4825_ (.A1(_4404_),
    .A2(_4405_),
    .ZN(_4406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4826_ (.A1(\as2650.alu_op[0] ),
    .A2(_4261_),
    .ZN(_4407_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4827_ (.I(_4407_),
    .Z(_4408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4828_ (.A1(_4210_),
    .A2(_4408_),
    .ZN(_4409_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4829_ (.A1(_4216_),
    .A2(_4232_),
    .ZN(_4410_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4830_ (.A1(_4372_),
    .A2(_4172_),
    .A3(_4410_),
    .ZN(_4411_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4831_ (.A1(_4406_),
    .A2(_4409_),
    .A3(_4411_),
    .ZN(_4412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4832_ (.A1(_4403_),
    .A2(_4412_),
    .ZN(_4413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4833_ (.I(_4413_),
    .Z(_4414_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4834_ (.A1(_4374_),
    .A2(_4384_),
    .B(_4402_),
    .C(_4414_),
    .ZN(_4415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4835_ (.I(_4230_),
    .Z(_4416_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4836_ (.A1(_4356_),
    .A2(_4371_),
    .B(_4415_),
    .C(_4416_),
    .ZN(_4417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4837_ (.A1(_4354_),
    .A2(_4355_),
    .B(_4417_),
    .ZN(_4418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4838_ (.A1(_4352_),
    .A2(_4418_),
    .ZN(_4419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4839_ (.I(_4182_),
    .Z(_4420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4840_ (.I(_4172_),
    .Z(_4421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4841_ (.A1(_4421_),
    .A2(_4207_),
    .ZN(_4422_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4842_ (.I(_4235_),
    .ZN(_4423_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4843_ (.A1(_4423_),
    .A2(_4267_),
    .ZN(_4424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4844_ (.I(_4424_),
    .Z(_4425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4845_ (.I(\as2650.addr_buff[7] ),
    .Z(_4426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4846_ (.I(_4426_),
    .Z(_4427_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4847_ (.A1(_4427_),
    .A2(_4245_),
    .ZN(_4428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4848_ (.A1(_4425_),
    .A2(_4428_),
    .ZN(_4429_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4849_ (.A1(_4420_),
    .A2(_4422_),
    .A3(_4429_),
    .ZN(_4430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4850_ (.I(_4430_),
    .Z(_4431_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4851_ (.I(\as2650.addr_buff[5] ),
    .ZN(_4432_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4852_ (.A1(\as2650.addr_buff[6] ),
    .A2(_4432_),
    .ZN(_4433_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4853_ (.I(\as2650.addr_buff[6] ),
    .ZN(_4434_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4854_ (.A1(_4434_),
    .A2(\as2650.addr_buff[5] ),
    .ZN(_4435_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4855_ (.A1(_4433_),
    .A2(_4435_),
    .ZN(_4436_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4856_ (.A1(_4398_),
    .A2(_4436_),
    .Z(_4437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4857_ (.I(_4437_),
    .Z(_4438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4858_ (.A1(_4431_),
    .A2(_4438_),
    .ZN(_4439_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4859_ (.A1(_4350_),
    .A2(_4419_),
    .A3(_4439_),
    .ZN(_4440_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4860_ (.I(_4113_),
    .Z(_4441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4861_ (.I(_4441_),
    .Z(_4442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4862_ (.I(_4423_),
    .Z(_4443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4863_ (.I(_4241_),
    .Z(_4444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4864_ (.A1(_4443_),
    .A2(_4444_),
    .ZN(_4445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4865_ (.I(_4260_),
    .Z(_4446_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4866_ (.I(_4446_),
    .Z(_4447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4867_ (.A1(_4271_),
    .A2(_4447_),
    .ZN(_4448_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4868_ (.A1(_4442_),
    .A2(_4257_),
    .A3(_4445_),
    .A4(_4448_),
    .ZN(_4449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4869_ (.I(_4397_),
    .Z(_4450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4870_ (.I(\as2650.idx_ctrl[1] ),
    .Z(_4451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4871_ (.I(\as2650.idx_ctrl[0] ),
    .Z(_4452_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4872_ (.I(_4452_),
    .ZN(_4453_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4873_ (.A1(_4451_),
    .A2(_4453_),
    .ZN(_4454_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4874_ (.I(_4451_),
    .ZN(_4455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4875_ (.A1(_4455_),
    .A2(_4452_),
    .ZN(_4456_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4876_ (.A1(_4454_),
    .A2(_4456_),
    .ZN(_4457_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4877_ (.A1(_4450_),
    .A2(_4457_),
    .Z(_4458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4878_ (.I(_4458_),
    .Z(_4459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4879_ (.A1(_4449_),
    .A2(_4459_),
    .ZN(_4460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4880_ (.A1(_4440_),
    .A2(_4460_),
    .ZN(_4461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4881_ (.A1(_4348_),
    .A2(_4461_),
    .ZN(_4462_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4882_ (.A1(_4290_),
    .A2(_4347_),
    .B(_4462_),
    .ZN(_4463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4883_ (.A1(_4118_),
    .A2(_4224_),
    .ZN(_4464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4884_ (.I(_4168_),
    .Z(_4465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4885_ (.I(_4465_),
    .Z(_4466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4886_ (.I(_4466_),
    .Z(_4467_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4887_ (.I(\as2650.psu[0] ),
    .Z(_4468_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4888_ (.I(_4468_),
    .ZN(_4469_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4889_ (.I(\as2650.psu[1] ),
    .ZN(_4470_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4890_ (.A1(_4469_),
    .A2(_4470_),
    .ZN(_4471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4891_ (.I(_4471_),
    .Z(_4472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4892_ (.I(_4472_),
    .Z(_4473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4893_ (.I(_4473_),
    .Z(_4474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4894_ (.I(_4471_),
    .Z(_4475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4895_ (.I(_4475_),
    .Z(_4476_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4896_ (.I(\as2650.psu[1] ),
    .Z(_4477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4897_ (.I(_4468_),
    .Z(_4478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4898_ (.A1(_4477_),
    .A2(\as2650.stack[5][8] ),
    .B1(\as2650.stack[4][8] ),
    .B2(_4478_),
    .ZN(_4479_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4899_ (.A1(_4476_),
    .A2(_4479_),
    .ZN(_4480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4900_ (.A1(\as2650.stack[6][8] ),
    .A2(_4474_),
    .B(_4480_),
    .ZN(_4481_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4901_ (.A1(\as2650.psu[0] ),
    .A2(\as2650.psu[1] ),
    .ZN(_4482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4902_ (.I(_4482_),
    .Z(_4483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4903_ (.I(_4483_),
    .Z(_4484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4904_ (.I(_4484_),
    .Z(_4485_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4905_ (.I(\as2650.psu[2] ),
    .ZN(_4486_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4906_ (.A1(_4486_),
    .A2(_4483_),
    .Z(_4487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4907_ (.I(_4487_),
    .Z(_4488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4908_ (.I(_4488_),
    .Z(_4489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4909_ (.I(_4489_),
    .Z(_4490_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4910_ (.A1(\as2650.stack[7][8] ),
    .A2(_4485_),
    .B(_4490_),
    .ZN(_4491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4911_ (.A1(_4477_),
    .A2(\as2650.stack[1][8] ),
    .B1(\as2650.stack[0][8] ),
    .B2(_4478_),
    .ZN(_4492_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4912_ (.A1(_4474_),
    .A2(_4492_),
    .Z(_4493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4913_ (.I(\as2650.psu[2] ),
    .Z(_4494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4914_ (.I(_4494_),
    .Z(_4495_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4915_ (.A1(\as2650.psu[2] ),
    .A2(_4482_),
    .Z(_4496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4916_ (.I(_4496_),
    .Z(_4497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4917_ (.I(_4497_),
    .Z(_4498_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4918_ (.I(_4498_),
    .Z(_4499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4919_ (.A1(_4495_),
    .A2(\as2650.stack[3][8] ),
    .B1(\as2650.stack[2][8] ),
    .B2(_4474_),
    .C(_4499_),
    .ZN(_4500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4920_ (.A1(_4481_),
    .A2(_4491_),
    .B1(_4493_),
    .B2(_4500_),
    .ZN(_4501_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4921_ (.A1(_4464_),
    .A2(_4467_),
    .A3(_4501_),
    .ZN(_4502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4922_ (.I(_4354_),
    .Z(_4503_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4923_ (.A1(_4135_),
    .A2(_4217_),
    .A3(_4294_),
    .ZN(_4504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4924_ (.A1(_4132_),
    .A2(_4177_),
    .ZN(_4505_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4925_ (.A1(_4504_),
    .A2(_4505_),
    .ZN(_4506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4926_ (.I(_4506_),
    .Z(_4507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4927_ (.I(_4507_),
    .Z(_4508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4928_ (.I(_4508_),
    .Z(_4509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4929_ (.I(_4509_),
    .Z(_4510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4930_ (.A1(_4198_),
    .A2(_4312_),
    .ZN(_4511_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4931_ (.I(_4511_),
    .ZN(_4512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4932_ (.A1(_4309_),
    .A2(_4512_),
    .ZN(_4513_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4933_ (.A1(_4513_),
    .A2(_4505_),
    .ZN(_4514_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4934_ (.A1(_4169_),
    .A2(_4514_),
    .ZN(_4515_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4935_ (.A1(_4464_),
    .A2(_4515_),
    .ZN(_4516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4936_ (.I(_4516_),
    .Z(_4517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4937_ (.A1(_4503_),
    .A2(_4510_),
    .B(_4517_),
    .ZN(_4518_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4938_ (.A1(_4502_),
    .A2(_4518_),
    .ZN(_4519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4939_ (.A1(_4288_),
    .A2(_4463_),
    .B(_4519_),
    .C(_4286_),
    .ZN(_4520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4940_ (.A1(_4107_),
    .A2(_4287_),
    .B(_4520_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4941_ (.I(\as2650.r123[0][1] ),
    .ZN(_4521_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4942_ (.A1(_4377_),
    .A2(_4381_),
    .Z(_4522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4943_ (.A1(\as2650.holding_reg[1] ),
    .A2(_4319_),
    .ZN(_4523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4944_ (.A1(_4319_),
    .A2(_4522_),
    .B(_4523_),
    .ZN(_4524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4945_ (.I(_4524_),
    .Z(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4946_ (.A1(_4273_),
    .A2(_4377_),
    .A3(_4381_),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4947_ (.I(_4379_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4948_ (.A1(_0286_),
    .A2(_4273_),
    .B(_4319_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4949_ (.A1(\as2650.holding_reg[1] ),
    .A2(_4129_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4950_ (.A1(_0285_),
    .A2(_0287_),
    .B(_0288_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4951_ (.A1(_0284_),
    .A2(_0289_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4952_ (.I(_0290_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4953_ (.A1(_4315_),
    .A2(_4329_),
    .B(_4339_),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4954_ (.I(_4154_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4955_ (.I(_0293_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4956_ (.A1(_0294_),
    .A2(_4293_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4957_ (.A1(_0291_),
    .A2(_0292_),
    .B(_0295_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4958_ (.A1(_0291_),
    .A2(_0292_),
    .B(_0296_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4959_ (.I(_0289_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4960_ (.A1(_4524_),
    .A2(_0298_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4961_ (.I0(_4322_),
    .I1(_4397_),
    .S(_4129_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4962_ (.A1(_0300_),
    .A2(_4327_),
    .A3(_4328_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4963_ (.A1(_0300_),
    .A2(_4321_),
    .A3(_4324_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4964_ (.A1(_4336_),
    .A2(_0301_),
    .B(_0302_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4965_ (.A1(_0299_),
    .A2(_0303_),
    .B(_4333_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4966_ (.A1(_0299_),
    .A2(_0303_),
    .B(_0304_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4967_ (.I(_4338_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4968_ (.A1(_0284_),
    .A2(_0298_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4969_ (.A1(_4310_),
    .A2(_0307_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4970_ (.I(_4218_),
    .Z(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4971_ (.A1(_0284_),
    .A2(_0298_),
    .B(_0308_),
    .C(_0309_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4972_ (.I(_4296_),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4973_ (.A1(_0306_),
    .A2(_0291_),
    .B(_0310_),
    .C(_0311_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _4974_ (.A1(_0297_),
    .A2(_0305_),
    .A3(_0312_),
    .B1(_0284_),
    .B2(_4298_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4975_ (.I(_4349_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4976_ (.I(_4305_),
    .Z(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4977_ (.I(_4522_),
    .Z(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4978_ (.A1(_4451_),
    .A2(_4453_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4979_ (.A1(_4450_),
    .A2(_4454_),
    .B(_0317_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4980_ (.A1(_0315_),
    .A2(_0316_),
    .A3(_0318_),
    .Z(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4981_ (.I(_0319_),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4982_ (.I(_4289_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4983_ (.A1(_0314_),
    .A2(_0320_),
    .B(_0321_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4984_ (.I(_4430_),
    .Z(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4985_ (.I(_4433_),
    .Z(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4986_ (.A1(_4243_),
    .A2(_4432_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4987_ (.A1(_0315_),
    .A2(_0324_),
    .B(_0325_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4988_ (.A1(_0315_),
    .A2(_4522_),
    .A3(_0326_),
    .Z(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4989_ (.I(_0327_),
    .Z(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4990_ (.I(_4379_),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4991_ (.I(_0329_),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4992_ (.I(_0330_),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4993_ (.I(_4406_),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4994_ (.I(_0332_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4995_ (.A1(_4217_),
    .A2(_4228_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4996_ (.A1(_4131_),
    .A2(_0334_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4997_ (.A1(_0333_),
    .A2(_4422_),
    .A3(_0335_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4998_ (.I(_0336_),
    .Z(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4999_ (.I(_4385_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5000_ (.I(_4375_),
    .Z(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5001_ (.I0(\as2650.r123[2][2] ),
    .I1(\as2650.r123_2[2][2] ),
    .S(_0339_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5002_ (.A1(_4361_),
    .A2(_0340_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5003_ (.I(\as2650.r0[2] ),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5004_ (.I(_0342_),
    .Z(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5005_ (.I0(\as2650.r123[1][2] ),
    .I1(\as2650.r123[0][2] ),
    .I2(\as2650.r123_2[1][2] ),
    .I3(\as2650.r123_2[0][2] ),
    .S0(_4366_),
    .S1(_0339_),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _5006_ (.A1(_0343_),
    .A2(_4175_),
    .B1(_4365_),
    .B2(_0344_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5007_ (.A1(_0341_),
    .A2(_0345_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5008_ (.I(_0346_),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5009_ (.I(_0347_),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5010_ (.I(net7),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5011_ (.I(_0349_),
    .Z(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5012_ (.I(_0350_),
    .Z(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5013_ (.I(_0351_),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5014_ (.I(_0352_),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5015_ (.I(_4395_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5016_ (.A1(\as2650.ins_reg[4] ),
    .A2(_4407_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5017_ (.I(_4450_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5018_ (.I(_4306_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5019_ (.A1(\as2650.ins_reg[4] ),
    .A2(_4262_),
    .A3(_0357_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5020_ (.A1(_0355_),
    .A2(_0356_),
    .B(_0358_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5021_ (.A1(_4384_),
    .A2(_0359_),
    .Z(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5022_ (.I(_0360_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5023_ (.A1(_0354_),
    .A2(_0361_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5024_ (.I(_4373_),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5025_ (.A1(_0353_),
    .A2(_0354_),
    .B(_0362_),
    .C(_0363_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5026_ (.I(_4414_),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5027_ (.A1(_0338_),
    .A2(_0348_),
    .B(_0364_),
    .C(_0365_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5028_ (.I(_0357_),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5029_ (.I(_0367_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5030_ (.I(_0336_),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5031_ (.A1(_4215_),
    .A2(_0368_),
    .B(_0369_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5032_ (.A1(_0331_),
    .A2(_0337_),
    .B1(_0366_),
    .B2(_0370_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5033_ (.A1(_0323_),
    .A2(_0371_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5034_ (.A1(_0323_),
    .A2(_0328_),
    .B(_0372_),
    .C(_4449_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5035_ (.A1(_4348_),
    .A2(_0313_),
    .B1(_0322_),
    .B2(_0373_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5036_ (.I(_4509_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5037_ (.A1(_4468_),
    .A2(\as2650.psu[1] ),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5038_ (.I(_0376_),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5039_ (.I(_4469_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5040_ (.I(_4470_),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5041_ (.A1(_0378_),
    .A2(_0379_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5042_ (.A1(_0377_),
    .A2(_0380_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5043_ (.I(_0381_),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5044_ (.I(_0378_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5045_ (.I(_0383_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5046_ (.I(_0379_),
    .Z(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5047_ (.I(_0385_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5048_ (.I(_0386_),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5049_ (.A1(_0384_),
    .A2(\as2650.stack[5][9] ),
    .B1(\as2650.stack[4][9] ),
    .B2(_0387_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5050_ (.A1(\as2650.stack[6][9] ),
    .A2(_4475_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5051_ (.A1(_0382_),
    .A2(_0388_),
    .B(_0389_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5052_ (.A1(\as2650.stack[7][9] ),
    .A2(_4484_),
    .B(_4489_),
    .C(_0390_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5053_ (.I(_4483_),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5054_ (.I(_0386_),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5055_ (.A1(_0384_),
    .A2(\as2650.stack[1][9] ),
    .B1(\as2650.stack[0][9] ),
    .B2(_0393_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5056_ (.A1(\as2650.stack[2][9] ),
    .A2(_4473_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5057_ (.A1(_0382_),
    .A2(_0394_),
    .B(_0395_),
    .C(_4489_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5058_ (.A1(\as2650.stack[3][9] ),
    .A2(_0392_),
    .B(_0396_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5059_ (.A1(_0391_),
    .A2(_0397_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5060_ (.A1(_0331_),
    .A2(_4510_),
    .B(_4517_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5061_ (.A1(_0375_),
    .A2(_0398_),
    .B(_0399_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5062_ (.I(_4285_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5063_ (.A1(_4288_),
    .A2(_0374_),
    .B(_0400_),
    .C(_0401_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5064_ (.A1(_4521_),
    .A2(_4287_),
    .B(_0402_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5065_ (.I(\as2650.r123[0][2] ),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5066_ (.I(_4236_),
    .Z(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5067_ (.A1(_0404_),
    .A2(_4404_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5068_ (.A1(_0405_),
    .A2(_4253_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5069_ (.A1(_4190_),
    .A2(_0406_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5070_ (.I(_0407_),
    .Z(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5071_ (.I(_0408_),
    .Z(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5072_ (.A1(_4442_),
    .A2(_4272_),
    .A3(_4264_),
    .A4(_0409_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5073_ (.A1(\as2650.holding_reg[2] ),
    .A2(_4320_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5074_ (.A1(_4161_),
    .A2(_0346_),
    .B(_0411_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5075_ (.A1(_4274_),
    .A2(_0341_),
    .A3(_0345_),
    .Z(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5076_ (.I(_0343_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5077_ (.A1(_0414_),
    .A2(_4275_),
    .B(_4320_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5078_ (.A1(\as2650.holding_reg[2] ),
    .A2(_4323_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5079_ (.A1(_0413_),
    .A2(_0415_),
    .B(_0416_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5080_ (.A1(_0412_),
    .A2(_0417_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5081_ (.A1(_0412_),
    .A2(_0417_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5082_ (.A1(_0418_),
    .A2(_0419_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5083_ (.I(_0420_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5084_ (.I(_4161_),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5085_ (.A1(_0422_),
    .A2(_0316_),
    .B(_4523_),
    .C(_0298_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5086_ (.A1(_0299_),
    .A2(_0303_),
    .B(_0423_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5087_ (.A1(_0421_),
    .A2(_0424_),
    .B(_4333_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5088_ (.A1(_0421_),
    .A2(_0424_),
    .B(_0425_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5089_ (.A1(_0290_),
    .A2(_0292_),
    .B(_0307_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5090_ (.A1(_0420_),
    .A2(_0427_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5091_ (.A1(_4313_),
    .A2(_0428_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5092_ (.A1(_4311_),
    .A2(_0309_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5093_ (.I(_4342_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5094_ (.I(_0418_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5095_ (.A1(_4292_),
    .A2(_4293_),
    .A3(_4295_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5096_ (.A1(_0431_),
    .A2(_0432_),
    .B(_0433_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _5097_ (.A1(_0430_),
    .A2(_0419_),
    .B1(_0421_),
    .B2(_4338_),
    .C(_0434_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5098_ (.I(_4297_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _5099_ (.A1(_0426_),
    .A2(_0429_),
    .A3(_0435_),
    .B1(_0412_),
    .B2(_0436_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5100_ (.I(_0414_),
    .Z(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5101_ (.I(_0438_),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5102_ (.I(_4356_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5103_ (.I(_0316_),
    .Z(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5104_ (.I(\as2650.r0[3] ),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5105_ (.I(_0442_),
    .Z(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5106_ (.I(_0443_),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5107_ (.A1(_0444_),
    .A2(_4176_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5108_ (.I0(\as2650.r123[2][3] ),
    .I1(\as2650.r123_2[2][3] ),
    .S(_0339_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5109_ (.A1(_4361_),
    .A2(_0446_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5110_ (.I0(\as2650.r123[1][3] ),
    .I1(\as2650.r123[0][3] ),
    .I2(\as2650.r123_2[1][3] ),
    .I3(\as2650.r123_2[0][3] ),
    .S0(_4366_),
    .S1(_4111_),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5111_ (.A1(_4365_),
    .A2(_0448_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5112_ (.A1(_0445_),
    .A2(_0447_),
    .A3(_0449_),
    .Z(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5113_ (.I(_0450_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5114_ (.I(_0451_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5115_ (.I(net8),
    .Z(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5116_ (.I(_0453_),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5117_ (.I(_0454_),
    .Z(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5118_ (.I(_0455_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5119_ (.I(_4395_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5120_ (.A1(_0341_),
    .A2(_0345_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5121_ (.I(_0458_),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5122_ (.A1(_4378_),
    .A2(_4382_),
    .B(_4397_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5123_ (.A1(_4384_),
    .A2(_0358_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5124_ (.A1(_4212_),
    .A2(_0460_),
    .B(_0461_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5125_ (.A1(_0459_),
    .A2(_0462_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5126_ (.A1(_4396_),
    .A2(_0463_),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5127_ (.A1(_0456_),
    .A2(_0457_),
    .B(_0464_),
    .C(_4385_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5128_ (.A1(_4374_),
    .A2(_0452_),
    .B(_0465_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5129_ (.A1(_4414_),
    .A2(_0466_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5130_ (.A1(_0440_),
    .A2(_0441_),
    .B(_0467_),
    .C(_4416_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5131_ (.A1(_0439_),
    .A2(_4355_),
    .B(_0468_),
    .C(_4351_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5132_ (.I(_4435_),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5133_ (.A1(_0315_),
    .A2(_4378_),
    .A3(_4382_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5134_ (.A1(_0458_),
    .A2(_0471_),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5135_ (.A1(_0346_),
    .A2(_0460_),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5136_ (.A1(_4436_),
    .A2(_0347_),
    .Z(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5137_ (.A1(_0470_),
    .A2(_0472_),
    .B1(_0473_),
    .B2(_0324_),
    .C(_0474_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5138_ (.I(_0475_),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5139_ (.A1(_4431_),
    .A2(_0476_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5140_ (.A1(_0314_),
    .A2(_0469_),
    .A3(_0477_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5141_ (.A1(_4456_),
    .A2(_0472_),
    .Z(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5142_ (.A1(_4455_),
    .A2(_4452_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5143_ (.A1(_0480_),
    .A2(_0317_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5144_ (.A1(_0458_),
    .A2(_0460_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5145_ (.I(_0480_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5146_ (.A1(_0481_),
    .A2(_0459_),
    .B1(_0482_),
    .B2(_0483_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5147_ (.A1(_0479_),
    .A2(_0484_),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5148_ (.A1(_4449_),
    .A2(_0485_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5149_ (.A1(_0478_),
    .A2(_0486_),
    .B(_0410_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5150_ (.A1(_0410_),
    .A2(_0437_),
    .B(_0487_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5151_ (.A1(\as2650.stack[7][10] ),
    .A2(_0392_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5152_ (.A1(_4499_),
    .A2(_0489_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5153_ (.I(_0381_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5154_ (.I(_0491_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5155_ (.I(_0378_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5156_ (.I(_0493_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5157_ (.I(_0494_),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5158_ (.I(_0387_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5159_ (.A1(_0495_),
    .A2(\as2650.stack[5][10] ),
    .B1(\as2650.stack[4][10] ),
    .B2(_0496_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5160_ (.A1(\as2650.stack[6][10] ),
    .A2(_4476_),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5161_ (.A1(_0492_),
    .A2(_0497_),
    .B(_0498_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5162_ (.A1(_0495_),
    .A2(\as2650.stack[1][10] ),
    .B1(\as2650.stack[0][10] ),
    .B2(_0496_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5163_ (.I(_4496_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5164_ (.I(_0501_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5165_ (.A1(_4494_),
    .A2(\as2650.stack[3][10] ),
    .B1(\as2650.stack[2][10] ),
    .B2(_4476_),
    .C(_0502_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5166_ (.A1(_0492_),
    .A2(_0500_),
    .B(_0503_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5167_ (.A1(_0490_),
    .A2(_0499_),
    .B(_0504_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5168_ (.I(_0439_),
    .Z(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5169_ (.I(_4508_),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5170_ (.A1(_0506_),
    .A2(_0507_),
    .B(_4516_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5171_ (.A1(_0375_),
    .A2(_0505_),
    .B(_0508_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5172_ (.A1(_4288_),
    .A2(_0488_),
    .B(_0509_),
    .C(_0401_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5173_ (.A1(_0403_),
    .A2(_4287_),
    .B(_0510_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5174_ (.I(\as2650.r123[0][3] ),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5175_ (.I(_4283_),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5176_ (.A1(\as2650.holding_reg[3] ),
    .A2(_4161_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5177_ (.A1(_0422_),
    .A2(_0450_),
    .B(_0513_),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5178_ (.I(\as2650.holding_reg[3] ),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5179_ (.A1(_0445_),
    .A2(_0447_),
    .A3(_0449_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5180_ (.I(_0516_),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5181_ (.A1(_4275_),
    .A2(_0517_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5182_ (.I(_0444_),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5183_ (.A1(_0519_),
    .A2(_4259_),
    .B(_4323_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5184_ (.A1(_0515_),
    .A2(_4130_),
    .B1(_0518_),
    .B2(_0520_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5185_ (.A1(_0514_),
    .A2(_0521_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5186_ (.A1(_0514_),
    .A2(_0521_),
    .Z(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5187_ (.A1(_0522_),
    .A2(_0523_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5188_ (.I(_0417_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5189_ (.A1(_0412_),
    .A2(_0525_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5190_ (.A1(_0420_),
    .A2(_0424_),
    .B(_0526_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5191_ (.A1(_0524_),
    .A2(_0527_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5192_ (.A1(_0524_),
    .A2(_0527_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5193_ (.A1(_4334_),
    .A2(_0529_),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5194_ (.I(_0522_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5195_ (.A1(_0531_),
    .A2(_0523_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5196_ (.I(_0419_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5197_ (.A1(_0432_),
    .A2(_0427_),
    .B(_0533_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5198_ (.A1(_0532_),
    .A2(_0534_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5199_ (.I(_0295_),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5200_ (.A1(_0294_),
    .A2(_4218_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5201_ (.A1(_0537_),
    .A2(_0531_),
    .B1(_0532_),
    .B2(_4338_),
    .C(_4297_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5202_ (.A1(_4341_),
    .A2(_0523_),
    .B1(_0535_),
    .B2(_0536_),
    .C(_0538_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5203_ (.A1(_0528_),
    .A2(_0530_),
    .B(_0539_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5204_ (.A1(_0436_),
    .A2(_0514_),
    .B(_0540_),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5205_ (.I(_4349_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5206_ (.I(_0519_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5207_ (.I(\as2650.r0[4] ),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5208_ (.I(_0544_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5209_ (.A1(_0545_),
    .A2(_4175_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5210_ (.I0(\as2650.r123[2][4] ),
    .I1(\as2650.r123_2[2][4] ),
    .S(_4301_),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5211_ (.A1(_4300_),
    .A2(_0547_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5212_ (.I0(\as2650.r123[1][4] ),
    .I1(\as2650.r123[0][4] ),
    .I2(\as2650.r123_2[1][4] ),
    .I3(\as2650.r123_2[0][4] ),
    .S0(_4146_),
    .S1(_0339_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5213_ (.A1(_4303_),
    .A2(_0549_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5214_ (.A1(_0546_),
    .A2(_0548_),
    .A3(_0550_),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5215_ (.I(_0551_),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5216_ (.I(_0552_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5217_ (.I(net9),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5218_ (.I(_0554_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5219_ (.I(_0555_),
    .Z(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5220_ (.I(_0517_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _5221_ (.A1(_4378_),
    .A2(_4382_),
    .B1(_0341_),
    .B2(_0345_),
    .C(_4305_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5222_ (.A1(_0347_),
    .A2(_0461_),
    .B1(_0558_),
    .B2(_4212_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5223_ (.A1(_0557_),
    .A2(_0559_),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5224_ (.A1(_4396_),
    .A2(_0560_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5225_ (.A1(_0556_),
    .A2(_0457_),
    .B(_0561_),
    .C(_4374_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5226_ (.A1(_0363_),
    .A2(_0553_),
    .B(_0562_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5227_ (.A1(_0365_),
    .A2(_0563_),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5228_ (.A1(_0440_),
    .A2(_0348_),
    .B(_0564_),
    .C(_4416_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5229_ (.A1(_0543_),
    .A2(_4355_),
    .B(_0565_),
    .C(_4352_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5230_ (.I(_4436_),
    .Z(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _5231_ (.A1(_0357_),
    .A2(_0316_),
    .A3(_0346_),
    .A4(_0450_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5232_ (.A1(_0459_),
    .A2(_0471_),
    .B(_0557_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5233_ (.A1(_0568_),
    .A2(_0569_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5234_ (.A1(_4434_),
    .A2(_4244_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5235_ (.A1(_0558_),
    .A2(_0517_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5236_ (.A1(_0571_),
    .A2(_0572_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _5237_ (.A1(_0567_),
    .A2(_0451_),
    .B1(_0570_),
    .B2(_0470_),
    .C(_0573_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5238_ (.I(_0574_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5239_ (.A1(_4431_),
    .A2(_0575_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5240_ (.A1(_0566_),
    .A2(_0576_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5241_ (.I(_4456_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5242_ (.A1(_0578_),
    .A2(_0570_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5243_ (.A1(_0481_),
    .A2(_0557_),
    .B1(_0572_),
    .B2(_0483_),
    .C(_0579_),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5244_ (.A1(_4350_),
    .A2(_0580_),
    .B(_4289_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5245_ (.A1(_0542_),
    .A2(_0577_),
    .B(_0581_),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5246_ (.A1(_0410_),
    .A2(_0541_),
    .B(_0582_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5247_ (.I(_0381_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5248_ (.I(_0494_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5249_ (.I(_0387_),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5250_ (.A1(_0585_),
    .A2(\as2650.stack[5][11] ),
    .B1(\as2650.stack[4][11] ),
    .B2(_0586_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5251_ (.I(_4475_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5252_ (.A1(\as2650.stack[6][11] ),
    .A2(_0588_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5253_ (.A1(_0584_),
    .A2(_0587_),
    .B(_0589_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5254_ (.A1(\as2650.stack[7][11] ),
    .A2(_4485_),
    .B(_4490_),
    .C(_0590_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5255_ (.I(_0384_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5256_ (.A1(_0592_),
    .A2(\as2650.stack[1][11] ),
    .B1(\as2650.stack[0][11] ),
    .B2(_0586_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5257_ (.A1(\as2650.stack[2][11] ),
    .A2(_4476_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5258_ (.A1(_0584_),
    .A2(_0593_),
    .B(_0594_),
    .C(_4489_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5259_ (.A1(\as2650.stack[3][11] ),
    .A2(_4485_),
    .B(_0595_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5260_ (.A1(_0591_),
    .A2(_0596_),
    .Z(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5261_ (.I(_0543_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5262_ (.A1(_0598_),
    .A2(_0507_),
    .B(_4516_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5263_ (.A1(_0375_),
    .A2(_0597_),
    .B(_0599_),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5264_ (.A1(_0512_),
    .A2(_0583_),
    .B(_0600_),
    .C(_0401_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5265_ (.A1(_0511_),
    .A2(_4287_),
    .B(_0601_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5266_ (.I(\as2650.r123[0][4] ),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5267_ (.I(_4286_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5268_ (.A1(_0432_),
    .A2(_0427_),
    .B(_0523_),
    .C(_0533_),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5269_ (.A1(\as2650.holding_reg[4] ),
    .A2(_0422_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5270_ (.A1(_4162_),
    .A2(_0551_),
    .B(_0605_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5271_ (.I(\as2650.holding_reg[4] ),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5272_ (.A1(_0546_),
    .A2(_0548_),
    .A3(_0550_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5273_ (.I(_0608_),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5274_ (.A1(_4275_),
    .A2(_0609_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5275_ (.I(_0545_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5276_ (.I(_0611_),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5277_ (.A1(_0612_),
    .A2(_4259_),
    .B(_4323_),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5278_ (.A1(_0607_),
    .A2(_4130_),
    .B1(_0610_),
    .B2(_0613_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5279_ (.I(_0614_),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5280_ (.A1(_0606_),
    .A2(_0615_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5281_ (.A1(_0531_),
    .A2(_0604_),
    .B(_0616_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5282_ (.A1(_0531_),
    .A2(_0616_),
    .A3(_0604_),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5283_ (.A1(_0536_),
    .A2(_0617_),
    .A3(_0618_),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5284_ (.A1(_0294_),
    .A2(_4312_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5285_ (.I(_0616_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5286_ (.I(_0514_),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5287_ (.A1(_0622_),
    .A2(_0521_),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5288_ (.A1(_0524_),
    .A2(_0527_),
    .B(_0623_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5289_ (.A1(_0621_),
    .A2(_0624_),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5290_ (.A1(_0616_),
    .A2(_0624_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5291_ (.A1(_0620_),
    .A2(_0625_),
    .A3(_0626_),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5292_ (.I(_0606_),
    .Z(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5293_ (.A1(_0628_),
    .A2(_0614_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5294_ (.A1(_4310_),
    .A2(_0629_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5295_ (.A1(_0628_),
    .A2(_0614_),
    .B(_0630_),
    .C(_0309_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5296_ (.A1(_0306_),
    .A2(_0621_),
    .B(_0631_),
    .C(_0311_),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _5297_ (.A1(_0619_),
    .A2(_0627_),
    .A3(_0632_),
    .B1(_0628_),
    .B2(_0436_),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5298_ (.I(_0633_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5299_ (.I(_4457_),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5300_ (.A1(_0558_),
    .A2(_0517_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5301_ (.A1(_0609_),
    .A2(_0636_),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5302_ (.I(_0609_),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5303_ (.A1(_4383_),
    .A2(_0458_),
    .A3(_0516_),
    .A4(_0608_),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5304_ (.I(_0639_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5305_ (.A1(_0638_),
    .A2(_0568_),
    .B1(_0640_),
    .B2(_0367_),
    .C(_0317_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5306_ (.A1(_0635_),
    .A2(_0552_),
    .B1(_0637_),
    .B2(_4454_),
    .C(_0641_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5307_ (.I(_0642_),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5308_ (.I(_0612_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5309_ (.I(\as2650.r123[0][5] ),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5310_ (.A1(_4375_),
    .A2(\as2650.r123_2[0][5] ),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5311_ (.A1(_4301_),
    .A2(_0645_),
    .B(_0646_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5312_ (.I(_0647_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5313_ (.I(_0648_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5314_ (.I(\as2650.r0[5] ),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5315_ (.I(_0650_),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5316_ (.I0(\as2650.r123[2][5] ),
    .I1(\as2650.r123_2[2][5] ),
    .S(_4111_),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5317_ (.A1(_4361_),
    .A2(_0652_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5318_ (.A1(_0651_),
    .A2(_4165_),
    .B(_0653_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5319_ (.A1(_4147_),
    .A2(_4149_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5320_ (.A1(_4403_),
    .A2(\as2650.r123_2[1][5] ),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5321_ (.I(_4110_),
    .Z(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5322_ (.A1(_0657_),
    .A2(\as2650.r123[1][5] ),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5323_ (.A1(_0655_),
    .A2(_0656_),
    .A3(_0658_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _5324_ (.A1(_4151_),
    .A2(_0649_),
    .B(_0654_),
    .C(_0659_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5325_ (.I(_0660_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5326_ (.I(_0661_),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5327_ (.I(_0662_),
    .Z(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5328_ (.I(_0663_),
    .Z(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5329_ (.I(_0664_),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5330_ (.A1(_4422_),
    .A2(_4203_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5331_ (.A1(_4136_),
    .A2(_4262_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5332_ (.A1(_4450_),
    .A2(_0639_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5333_ (.A1(_0558_),
    .A2(_0516_),
    .A3(_0609_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5334_ (.I(_0355_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5335_ (.A1(_0670_),
    .A2(_0636_),
    .B(_0552_),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5336_ (.A1(_0667_),
    .A2(_0568_),
    .B1(_0669_),
    .B2(_0670_),
    .C(_0671_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5337_ (.A1(_0667_),
    .A2(_0668_),
    .B(_0672_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5338_ (.I(net10),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5339_ (.I(_0674_),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5340_ (.I(_0675_),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5341_ (.I(_0676_),
    .Z(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5342_ (.A1(_0677_),
    .A2(_0457_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5343_ (.A1(_0666_),
    .A2(_0673_),
    .B(_0678_),
    .C(_0338_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5344_ (.A1(_0338_),
    .A2(_0665_),
    .B(_0679_),
    .C(_0365_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5345_ (.I(_0452_),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5346_ (.A1(_4215_),
    .A2(_0681_),
    .B(_0369_),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5347_ (.A1(_0644_),
    .A2(_0337_),
    .B1(_0680_),
    .B2(_0682_),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5348_ (.A1(_0638_),
    .A2(_0568_),
    .B1(_0640_),
    .B2(_0356_),
    .C(_0325_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5349_ (.A1(_0567_),
    .A2(_0552_),
    .B1(_0637_),
    .B2(_0324_),
    .C(_0684_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5350_ (.I(_0685_),
    .Z(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5351_ (.A1(_4431_),
    .A2(_0686_),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5352_ (.A1(_0323_),
    .A2(_0683_),
    .B(_0687_),
    .C(_4350_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5353_ (.A1(_0542_),
    .A2(_0643_),
    .B(_0688_),
    .C(_0321_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5354_ (.A1(_4348_),
    .A2(_0634_),
    .B(_0689_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5355_ (.I(_4367_),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5356_ (.I(_4164_),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5357_ (.A1(_0691_),
    .A2(_0692_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5358_ (.A1(_4227_),
    .A2(_4513_),
    .A3(_0693_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5359_ (.A1(_0694_),
    .A2(_4506_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5360_ (.A1(_4145_),
    .A2(_4167_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5361_ (.A1(_0695_),
    .A2(_0696_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5362_ (.A1(_4127_),
    .A2(_0697_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5363_ (.I(_0644_),
    .Z(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5364_ (.A1(_0699_),
    .A2(_4509_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5365_ (.A1(_0592_),
    .A2(\as2650.stack[1][12] ),
    .B1(\as2650.stack[0][12] ),
    .B2(_0496_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5366_ (.A1(_0392_),
    .A2(_0701_),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5367_ (.A1(_4495_),
    .A2(\as2650.stack[3][12] ),
    .B1(\as2650.stack[2][12] ),
    .B2(_4474_),
    .C(_0502_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5368_ (.A1(_0585_),
    .A2(\as2650.stack[5][12] ),
    .B1(\as2650.stack[4][12] ),
    .B2(_0393_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5369_ (.A1(\as2650.stack[6][12] ),
    .A2(_4473_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5370_ (.A1(_0491_),
    .A2(_0704_),
    .B(_0705_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5371_ (.A1(\as2650.stack[7][12] ),
    .A2(_4485_),
    .B(_4490_),
    .C(_0706_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5372_ (.A1(_0702_),
    .A2(_0703_),
    .B(_0707_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5373_ (.A1(_4467_),
    .A2(_0708_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5374_ (.A1(_0698_),
    .A2(_0700_),
    .A3(_0709_),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5375_ (.A1(_0512_),
    .A2(_0690_),
    .B(_0710_),
    .C(_0401_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5376_ (.A1(_0602_),
    .A2(_0603_),
    .B(_0711_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5377_ (.I(_0422_),
    .Z(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5378_ (.A1(\as2650.holding_reg[5] ),
    .A2(_0712_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5379_ (.A1(_0712_),
    .A2(_0662_),
    .B(_0713_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5380_ (.I(_0650_),
    .Z(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5381_ (.I(_0715_),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5382_ (.A1(_4276_),
    .A2(_0661_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5383_ (.A1(_0716_),
    .A2(_4276_),
    .B(_0717_),
    .C(_4162_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5384_ (.A1(\as2650.holding_reg[5] ),
    .A2(_4130_),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5385_ (.A1(_0718_),
    .A2(_0719_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5386_ (.A1(_0714_),
    .A2(_0720_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5387_ (.I(_0721_),
    .Z(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5388_ (.A1(_0628_),
    .A2(_0615_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5389_ (.A1(_0626_),
    .A2(_0722_),
    .A3(_0723_),
    .Z(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5390_ (.A1(_0626_),
    .A2(_0723_),
    .B(_0721_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5391_ (.A1(_4334_),
    .A2(_0724_),
    .A3(_0725_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5392_ (.A1(_0629_),
    .A2(_0618_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5393_ (.A1(_0722_),
    .A2(_0727_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5394_ (.I(_0714_),
    .Z(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5395_ (.A1(_0729_),
    .A2(_0720_),
    .Z(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5396_ (.A1(_0729_),
    .A2(_0720_),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5397_ (.A1(_4341_),
    .A2(_0730_),
    .B1(_0731_),
    .B2(_0431_),
    .C(_0433_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5398_ (.A1(_0306_),
    .A2(_0722_),
    .B(_0732_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5399_ (.A1(_0536_),
    .A2(_0728_),
    .B(_0733_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5400_ (.A1(_0436_),
    .A2(_0729_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5401_ (.A1(_0726_),
    .A2(_0734_),
    .B(_0735_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5402_ (.A1(_0668_),
    .A2(_0660_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5403_ (.A1(_0669_),
    .A2(_0660_),
    .Z(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5404_ (.A1(_0571_),
    .A2(_0738_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5405_ (.A1(_4436_),
    .A2(_0662_),
    .B1(_0737_),
    .B2(_0470_),
    .C(_0739_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5406_ (.I(_0740_),
    .Z(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5407_ (.I(_0638_),
    .Z(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5408_ (.I(\as2650.r0[6] ),
    .Z(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5409_ (.I(_0743_),
    .Z(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5410_ (.I(_0744_),
    .Z(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5411_ (.A1(_0745_),
    .A2(_4176_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5412_ (.I0(\as2650.r123[2][6] ),
    .I1(\as2650.r123_2[2][6] ),
    .S(_0657_),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5413_ (.A1(_4362_),
    .A2(_0747_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5414_ (.I0(\as2650.r123[1][6] ),
    .I1(\as2650.r123[0][6] ),
    .I2(\as2650.r123_2[1][6] ),
    .I3(\as2650.r123_2[0][6] ),
    .S0(_4366_),
    .S1(_4112_),
    .Z(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5415_ (.A1(_4365_),
    .A2(_0749_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5416_ (.A1(_0746_),
    .A2(_0748_),
    .A3(_0750_),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5417_ (.I(_0751_),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5418_ (.I(_0752_),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5419_ (.I(_0753_),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5420_ (.I(net1),
    .Z(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5421_ (.I(_0755_),
    .Z(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5422_ (.I(_0756_),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5423_ (.I(_0757_),
    .Z(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5424_ (.A1(_0670_),
    .A2(_0669_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5425_ (.A1(_4136_),
    .A2(_4263_),
    .A3(_0356_),
    .A4(_0640_),
    .Z(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5426_ (.A1(_0759_),
    .A2(_0760_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5427_ (.A1(_0663_),
    .A2(_0761_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5428_ (.A1(_4396_),
    .A2(_0762_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5429_ (.A1(_0758_),
    .A2(_0354_),
    .B(_0763_),
    .C(_4374_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5430_ (.A1(_0363_),
    .A2(_0754_),
    .B(_0764_),
    .C(_4414_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5431_ (.A1(_0440_),
    .A2(_0742_),
    .B(_0765_),
    .C(_4416_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5432_ (.A1(_0651_),
    .A2(_4355_),
    .B(_0766_),
    .C(_4351_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5433_ (.A1(_4352_),
    .A2(_0741_),
    .B(_0767_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5434_ (.A1(_0483_),
    .A2(_0738_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5435_ (.A1(_0635_),
    .A2(_0663_),
    .B1(_0737_),
    .B2(_0578_),
    .C(_0769_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5436_ (.I(_0770_),
    .Z(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5437_ (.A1(_4350_),
    .A2(_0771_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5438_ (.A1(_0314_),
    .A2(_0768_),
    .B(_0772_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5439_ (.I0(_0736_),
    .I1(_0773_),
    .S(_0321_),
    .Z(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5440_ (.A1(_0585_),
    .A2(\as2650.stack[5][13] ),
    .B1(\as2650.stack[4][13] ),
    .B2(_0393_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5441_ (.A1(\as2650.stack[6][13] ),
    .A2(_0588_),
    .B1(_4484_),
    .B2(\as2650.stack[7][13] ),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5442_ (.A1(_0491_),
    .A2(_0775_),
    .B(_0776_),
    .C(_0502_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5443_ (.A1(_0592_),
    .A2(\as2650.stack[1][13] ),
    .B1(\as2650.stack[0][13] ),
    .B2(_0586_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5444_ (.A1(\as2650.stack[2][13] ),
    .A2(_0588_),
    .B1(_4484_),
    .B2(\as2650.stack[3][13] ),
    .C(_0502_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5445_ (.A1(_0584_),
    .A2(_0778_),
    .B(_0779_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5446_ (.A1(_0777_),
    .A2(_0780_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5447_ (.I(_0716_),
    .Z(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5448_ (.I(_0782_),
    .Z(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5449_ (.I(_0783_),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5450_ (.A1(_0784_),
    .A2(_0507_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5451_ (.A1(_4510_),
    .A2(_0781_),
    .B(_0785_),
    .C(_0698_),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5452_ (.A1(_0512_),
    .A2(_0774_),
    .B(_0786_),
    .C(_4285_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5453_ (.A1(_0645_),
    .A2(_0603_),
    .B(_0787_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5454_ (.I(\as2650.r123[0][6] ),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5455_ (.A1(\as2650.holding_reg[6] ),
    .A2(_4162_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5456_ (.A1(_0712_),
    .A2(_0751_),
    .B(_0789_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5457_ (.A1(_0746_),
    .A2(_0748_),
    .A3(_0750_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5458_ (.I(_0791_),
    .Z(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5459_ (.I(_0745_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5460_ (.A1(_0793_),
    .A2(_4260_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5461_ (.A1(_4260_),
    .A2(_0792_),
    .B(_0794_),
    .C(_0712_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5462_ (.A1(\as2650.holding_reg[6] ),
    .A2(_4131_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5463_ (.A1(_0795_),
    .A2(_0796_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5464_ (.A1(_0790_),
    .A2(_0797_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5465_ (.I(_0790_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5466_ (.A1(_0799_),
    .A2(_0795_),
    .A3(_0796_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5467_ (.A1(_0798_),
    .A2(_0800_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5468_ (.I(_0801_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5469_ (.A1(_0731_),
    .A2(_0727_),
    .B(_0730_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5470_ (.A1(_0802_),
    .A2(_0803_),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5471_ (.A1(_4313_),
    .A2(_0804_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5472_ (.A1(_0718_),
    .A2(_0719_),
    .B(_0729_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5473_ (.I(_0806_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5474_ (.A1(_0725_),
    .A2(_0807_),
    .B(_0802_),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5475_ (.A1(_0725_),
    .A2(_0802_),
    .A3(_0807_),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5476_ (.A1(_0620_),
    .A2(_0808_),
    .A3(_0809_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5477_ (.A1(_4310_),
    .A2(_0798_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5478_ (.A1(_0309_),
    .A2(_0800_),
    .A3(_0811_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5479_ (.A1(_0306_),
    .A2(_0801_),
    .B(_0812_),
    .C(_0311_),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _5480_ (.A1(_0805_),
    .A2(_0810_),
    .A3(_0813_),
    .B1(_0790_),
    .B2(_4298_),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5481_ (.A1(_0357_),
    .A2(_0639_),
    .A3(_0661_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5482_ (.A1(_0815_),
    .A2(_0791_),
    .Z(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5483_ (.A1(_0669_),
    .A2(_0660_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5484_ (.A1(_0817_),
    .A2(_0791_),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5485_ (.A1(_0483_),
    .A2(_0818_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5486_ (.A1(_0635_),
    .A2(_0752_),
    .B1(_0816_),
    .B2(_0578_),
    .C(_0819_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5487_ (.I(_0820_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5488_ (.I(_0745_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5489_ (.I(_0822_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5490_ (.A1(_4360_),
    .A2(_4364_),
    .A3(_4369_),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5491_ (.I(_0824_),
    .Z(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5492_ (.I(_0825_),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5493_ (.I(_0826_),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5494_ (.I0(_0759_),
    .I1(_0760_),
    .S(_0662_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5495_ (.A1(_0792_),
    .A2(_0828_),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5496_ (.I(net2),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5497_ (.I(_0830_),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5498_ (.I(_0831_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5499_ (.I(_0832_),
    .Z(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5500_ (.A1(_0833_),
    .A2(_0457_),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5501_ (.A1(_0666_),
    .A2(_0829_),
    .B(_0834_),
    .C(_0363_),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5502_ (.A1(_0338_),
    .A2(_0827_),
    .B(_0835_),
    .C(_0365_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5503_ (.A1(_4215_),
    .A2(_0665_),
    .B(_0369_),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5504_ (.A1(_0823_),
    .A2(_0337_),
    .B1(_0836_),
    .B2(_0837_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5505_ (.A1(_0571_),
    .A2(_0818_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5506_ (.A1(_0567_),
    .A2(_0753_),
    .B1(_0816_),
    .B2(_0470_),
    .C(_0839_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5507_ (.I(_0840_),
    .Z(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5508_ (.A1(_4430_),
    .A2(_0841_),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5509_ (.A1(_0323_),
    .A2(_0838_),
    .B(_0842_),
    .C(_4349_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5510_ (.A1(_0542_),
    .A2(_0821_),
    .B(_0843_),
    .C(_0321_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5511_ (.A1(_4348_),
    .A2(_0814_),
    .B(_0844_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5512_ (.A1(\as2650.stack[7][14] ),
    .A2(_0392_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5513_ (.A1(_0384_),
    .A2(\as2650.stack[5][14] ),
    .B1(\as2650.stack[4][14] ),
    .B2(_0387_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5514_ (.A1(_0382_),
    .A2(_0847_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5515_ (.A1(\as2650.stack[6][14] ),
    .A2(_0588_),
    .B(_0848_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5516_ (.A1(_4499_),
    .A2(_0846_),
    .A3(_0849_),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5517_ (.A1(_0592_),
    .A2(\as2650.stack[1][14] ),
    .B1(\as2650.stack[0][14] ),
    .B2(_0586_),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5518_ (.A1(_4494_),
    .A2(\as2650.stack[3][14] ),
    .B1(\as2650.stack[2][14] ),
    .B2(_4473_),
    .C(_4498_),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5519_ (.A1(_0584_),
    .A2(_0851_),
    .B(_0852_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5520_ (.A1(_0850_),
    .A2(_0853_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5521_ (.A1(_0823_),
    .A2(_0507_),
    .B(_4516_),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5522_ (.A1(_0375_),
    .A2(_0854_),
    .B(_0855_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5523_ (.A1(_0512_),
    .A2(_0845_),
    .B(_0856_),
    .C(_4285_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5524_ (.A1(_0788_),
    .A2(_0603_),
    .B(_0857_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5525_ (.I(\as2650.r123[0][7] ),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5526_ (.I(_4359_),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5527_ (.I(_0859_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5528_ (.I(_0860_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5529_ (.I(_0861_),
    .Z(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5530_ (.A1(_0862_),
    .A2(_4467_),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5531_ (.A1(_4517_),
    .A2(_0863_),
    .B(_4286_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5532_ (.A1(\as2650.holding_reg[7] ),
    .A2(_4163_),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5533_ (.A1(_4226_),
    .A2(_0826_),
    .B(_0865_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5534_ (.A1(_4276_),
    .A2(_0825_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5535_ (.A1(_4359_),
    .A2(_4277_),
    .B(_0867_),
    .C(_4163_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5536_ (.A1(\as2650.holding_reg[7] ),
    .A2(_4131_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5537_ (.A1(_0868_),
    .A2(_0869_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5538_ (.A1(_0866_),
    .A2(_0870_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5539_ (.A1(_0866_),
    .A2(_0870_),
    .Z(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5540_ (.A1(_0871_),
    .A2(_0872_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5541_ (.A1(_0798_),
    .A2(_0803_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5542_ (.A1(_0800_),
    .A2(_0874_),
    .Z(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5543_ (.A1(_0873_),
    .A2(_0875_),
    .Z(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5544_ (.A1(_0799_),
    .A2(_0797_),
    .B(_0808_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5545_ (.A1(_0873_),
    .A2(_0877_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5546_ (.I(_0871_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5547_ (.A1(_4295_),
    .A2(_0873_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5548_ (.A1(_4341_),
    .A2(_0879_),
    .B1(_0872_),
    .B2(_0431_),
    .C(_0880_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5549_ (.A1(_4313_),
    .A2(_0876_),
    .B1(_0878_),
    .B2(_0620_),
    .C(_0881_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5550_ (.I0(_0866_),
    .I1(_0882_),
    .S(_0311_),
    .Z(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5551_ (.I(_0883_),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5552_ (.A1(_0817_),
    .A2(_0791_),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5553_ (.A1(_4370_),
    .A2(_0885_),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5554_ (.A1(_0356_),
    .A2(_0639_),
    .A3(_0661_),
    .A4(_0751_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5555_ (.A1(_0824_),
    .A2(_0887_),
    .Z(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5556_ (.A1(_0317_),
    .A2(_0888_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5557_ (.A1(_0825_),
    .A2(_0635_),
    .B1(_0886_),
    .B2(_4454_),
    .C(_0889_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5558_ (.I(_0890_),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5559_ (.A1(_0325_),
    .A2(_0888_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _5560_ (.A1(_0825_),
    .A2(_0567_),
    .B1(_0886_),
    .B2(_0324_),
    .C(_0892_),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5561_ (.I(_0893_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5562_ (.A1(_0667_),
    .A2(_0815_),
    .Z(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5563_ (.A1(_4212_),
    .A2(_0817_),
    .B(_0752_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5564_ (.A1(_0895_),
    .A2(_0752_),
    .B(_0896_),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5565_ (.A1(_4370_),
    .A2(_0897_),
    .Z(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5566_ (.A1(_0666_),
    .A2(_0898_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5567_ (.I(net3),
    .Z(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5568_ (.I(_0900_),
    .Z(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5569_ (.I(_0901_),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5570_ (.A1(_0902_),
    .A2(_0354_),
    .B(_4223_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5571_ (.A1(_4357_),
    .A2(_4398_),
    .B(_4336_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5572_ (.I(_0904_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5573_ (.A1(_0899_),
    .A2(_0903_),
    .B1(_0905_),
    .B2(_4223_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5574_ (.A1(_4356_),
    .A2(_0754_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5575_ (.A1(_0440_),
    .A2(_0906_),
    .B(_0907_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5576_ (.I(_0860_),
    .Z(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5577_ (.A1(_0909_),
    .A2(_0369_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5578_ (.A1(_0337_),
    .A2(_0908_),
    .B(_0910_),
    .C(_4351_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5579_ (.A1(_4352_),
    .A2(_0894_),
    .B(_0911_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5580_ (.A1(_0314_),
    .A2(_0912_),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5581_ (.A1(_0542_),
    .A2(_0891_),
    .B(_0913_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5582_ (.A1(_4290_),
    .A2(_0914_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5583_ (.A1(_4290_),
    .A2(_0884_),
    .B(_0915_),
    .C(_4288_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5584_ (.A1(_0858_),
    .A2(_0603_),
    .B1(_0864_),
    .B2(_0916_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5585_ (.I(_4477_),
    .Z(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5586_ (.I(_4486_),
    .Z(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5587_ (.I(_0918_),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5588_ (.A1(_0917_),
    .A2(_0919_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5589_ (.I(_4197_),
    .Z(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5590_ (.I(_0921_),
    .Z(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5591_ (.A1(_4512_),
    .A2(_4362_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5592_ (.A1(_4390_),
    .A2(_0923_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5593_ (.A1(_0922_),
    .A2(_0924_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5594_ (.I(_4404_),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5595_ (.I(_4189_),
    .Z(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _5596_ (.A1(_4238_),
    .A2(_0927_),
    .A3(_0404_),
    .A4(_4190_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5597_ (.A1(_0926_),
    .A2(_0928_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5598_ (.I(_0921_),
    .Z(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5599_ (.I(_4389_),
    .Z(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5600_ (.A1(_0930_),
    .A2(_0931_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5601_ (.I(net3),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5602_ (.A1(_0925_),
    .A2(_0929_),
    .B1(_0932_),
    .B2(_0933_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5603_ (.I(_4255_),
    .Z(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5604_ (.A1(_4426_),
    .A2(_0935_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5605_ (.A1(_0293_),
    .A2(_0925_),
    .B(_0936_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5606_ (.I(_4209_),
    .Z(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5607_ (.A1(_0938_),
    .A2(_0924_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5608_ (.A1(_4185_),
    .A2(_0939_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5609_ (.A1(_0293_),
    .A2(_4182_),
    .A3(_4261_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5610_ (.A1(_0934_),
    .A2(_0937_),
    .B(_0940_),
    .C(_0941_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5611_ (.I(_4192_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5612_ (.A1(_0943_),
    .A2(_0926_),
    .A3(_4123_),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5613_ (.I(_0944_),
    .Z(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5614_ (.A1(_4132_),
    .A2(_4151_),
    .A3(_4158_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5615_ (.A1(_0945_),
    .A2(_0946_),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5616_ (.I(_0925_),
    .Z(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5617_ (.A1(_4238_),
    .A2(_4189_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5618_ (.A1(_4252_),
    .A2(_0949_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5619_ (.A1(_4122_),
    .A2(_0950_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5620_ (.A1(_0293_),
    .A2(_0951_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5621_ (.A1(_0948_),
    .A2(_0952_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5622_ (.A1(_0942_),
    .A2(_0947_),
    .A3(_0953_),
    .B(_4421_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5623_ (.A1(_4478_),
    .A2(_0954_),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5624_ (.A1(_0920_),
    .A2(_0955_),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5625_ (.I(_0956_),
    .Z(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5626_ (.I(_0957_),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5627_ (.I0(\as2650.r123[0][0] ),
    .I1(\as2650.r123_2[0][0] ),
    .S(_4109_),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5628_ (.I(_0959_),
    .Z(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5629_ (.I(_0960_),
    .Z(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5630_ (.I(_0961_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5631_ (.I(_4421_),
    .Z(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5632_ (.A1(_0963_),
    .A2(_0947_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5633_ (.I(_0964_),
    .Z(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5634_ (.I(\as2650.pc[8] ),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5635_ (.I(_0966_),
    .Z(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5636_ (.I(_0967_),
    .Z(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5637_ (.I(_0944_),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5638_ (.I(_0969_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5639_ (.I(_0946_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5640_ (.I(_0971_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5641_ (.A1(_4270_),
    .A2(_0970_),
    .A3(_0972_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5642_ (.I(_0973_),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5643_ (.A1(_0968_),
    .A2(_0974_),
    .Z(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5644_ (.A1(_0962_),
    .A2(_0965_),
    .B(_0975_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5645_ (.I(_0976_),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5646_ (.I(_0957_),
    .Z(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5647_ (.A1(\as2650.stack[2][8] ),
    .A2(_0978_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5648_ (.A1(_0958_),
    .A2(_0977_),
    .B(_0979_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5649_ (.I0(\as2650.r123[0][1] ),
    .I1(\as2650.r123_2[0][1] ),
    .S(_4108_),
    .Z(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5650_ (.I(_0980_),
    .Z(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5651_ (.I(_0981_),
    .Z(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5652_ (.I(_0982_),
    .Z(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5653_ (.I(_0983_),
    .Z(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5654_ (.I(\as2650.pc[9] ),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5655_ (.I(_0985_),
    .Z(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5656_ (.I(_0964_),
    .Z(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5657_ (.A1(_0986_),
    .A2(_0987_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5658_ (.A1(_0984_),
    .A2(_0965_),
    .B(_0988_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5659_ (.I(_0989_),
    .Z(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5660_ (.I(_0956_),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5661_ (.A1(\as2650.stack[2][9] ),
    .A2(_0991_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5662_ (.A1(_0958_),
    .A2(_0990_),
    .B(_0992_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5663_ (.I0(\as2650.r123[0][2] ),
    .I1(\as2650.r123_2[0][2] ),
    .S(\as2650.psl[4] ),
    .Z(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5664_ (.I(_0993_),
    .Z(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5665_ (.I(_0994_),
    .Z(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5666_ (.I(_0995_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5667_ (.I(\as2650.pc[10] ),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5668_ (.I(_0997_),
    .Z(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5669_ (.A1(_0998_),
    .A2(_0987_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5670_ (.A1(_0996_),
    .A2(_0965_),
    .B(_0999_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5671_ (.I(_1000_),
    .Z(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5672_ (.A1(\as2650.stack[2][10] ),
    .A2(_0991_),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5673_ (.A1(_0958_),
    .A2(_1001_),
    .B(_1002_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5674_ (.A1(_0657_),
    .A2(\as2650.r123_2[0][3] ),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5675_ (.A1(_0657_),
    .A2(_0511_),
    .B(_1003_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5676_ (.I(_1004_),
    .Z(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5677_ (.I(_1005_),
    .Z(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5678_ (.I(_1006_),
    .Z(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5679_ (.I(\as2650.pc[11] ),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5680_ (.I(_0964_),
    .Z(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5681_ (.A1(_1008_),
    .A2(_1009_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5682_ (.A1(_1007_),
    .A2(_0965_),
    .B(_1010_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5683_ (.I(_1011_),
    .Z(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5684_ (.A1(\as2650.stack[2][11] ),
    .A2(_0991_),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5685_ (.A1(_0958_),
    .A2(_1012_),
    .B(_1013_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5686_ (.I0(\as2650.r123[0][4] ),
    .I1(\as2650.r123_2[0][4] ),
    .S(_4108_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5687_ (.I(_1014_),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5688_ (.I(_1015_),
    .Z(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5689_ (.I(\as2650.pc[12] ),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5690_ (.I(_1017_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5691_ (.A1(_1018_),
    .A2(_1009_),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5692_ (.A1(_1016_),
    .A2(_0987_),
    .B(_1019_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5693_ (.I(_1020_),
    .Z(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5694_ (.A1(\as2650.stack[2][12] ),
    .A2(_0991_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5695_ (.A1(_0978_),
    .A2(_1021_),
    .B(_1022_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5696_ (.I(_0649_),
    .Z(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5697_ (.I(_1023_),
    .Z(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5698_ (.I(\as2650.pc[13] ),
    .Z(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5699_ (.A1(_1025_),
    .A2(_0974_),
    .Z(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5700_ (.A1(_1024_),
    .A2(_0987_),
    .B(_1026_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5701_ (.I(_1027_),
    .Z(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5702_ (.A1(\as2650.stack[2][13] ),
    .A2(_0957_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5703_ (.A1(_0978_),
    .A2(_1028_),
    .B(_1029_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5704_ (.I(\as2650.pc[14] ),
    .Z(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5705_ (.I(_4270_),
    .Z(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5706_ (.A1(_0332_),
    .A2(_0946_),
    .Z(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5707_ (.I(_1032_),
    .Z(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5708_ (.A1(_1031_),
    .A2(_1033_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5709_ (.I(_1034_),
    .Z(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5710_ (.A1(_4109_),
    .A2(\as2650.r123_2[0][6] ),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5711_ (.A1(_4110_),
    .A2(_0788_),
    .B(_1036_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5712_ (.I(_1037_),
    .Z(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5713_ (.I(_1038_),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5714_ (.I(_1039_),
    .Z(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5715_ (.A1(_1031_),
    .A2(_1040_),
    .A3(_1033_),
    .Z(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5716_ (.A1(_1030_),
    .A2(_1035_),
    .B(_1041_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5717_ (.I(_1042_),
    .Z(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5718_ (.A1(\as2650.stack[2][14] ),
    .A2(_0957_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5719_ (.A1(_0978_),
    .A2(_1043_),
    .B(_1044_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5720_ (.I(_0393_),
    .Z(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5721_ (.I(_1045_),
    .Z(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5722_ (.I(_0919_),
    .Z(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5723_ (.I(_1047_),
    .Z(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5724_ (.A1(_0585_),
    .A2(_0954_),
    .Z(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5725_ (.I(_1049_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5726_ (.I(_1050_),
    .Z(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5727_ (.A1(_1046_),
    .A2(_1048_),
    .A3(_1051_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5728_ (.I(_1052_),
    .Z(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5729_ (.I(_4503_),
    .Z(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5730_ (.I(\as2650.pc[0] ),
    .Z(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5731_ (.I(_1055_),
    .Z(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5732_ (.I(_1056_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5733_ (.I(_1057_),
    .Z(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5734_ (.I(_0973_),
    .Z(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5735_ (.A1(_1058_),
    .A2(_1059_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5736_ (.A1(_1054_),
    .A2(_1035_),
    .B(_1060_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5737_ (.I(_1061_),
    .Z(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5738_ (.I(_1052_),
    .Z(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5739_ (.A1(\as2650.stack[1][0] ),
    .A2(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5740_ (.A1(_1053_),
    .A2(_1062_),
    .B(_1064_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5741_ (.I(_0331_),
    .Z(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5742_ (.I(\as2650.pc[1] ),
    .Z(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5743_ (.I(_1066_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5744_ (.I(_1067_),
    .Z(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5745_ (.A1(_1068_),
    .A2(_1059_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5746_ (.A1(_1065_),
    .A2(_1035_),
    .B(_1069_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5747_ (.I(_1070_),
    .Z(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5748_ (.A1(\as2650.stack[1][1] ),
    .A2(_1063_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5749_ (.A1(_1053_),
    .A2(_1071_),
    .B(_1072_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5750_ (.I(\as2650.pc[2] ),
    .Z(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5751_ (.I(_1073_),
    .Z(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5752_ (.I(_1074_),
    .Z(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5753_ (.I(_1075_),
    .Z(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5754_ (.A1(_1076_),
    .A2(_1009_),
    .Z(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5755_ (.A1(_0506_),
    .A2(_1035_),
    .B(_1077_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5756_ (.I(_1078_),
    .Z(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5757_ (.A1(\as2650.stack[1][2] ),
    .A2(_1063_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5758_ (.A1(_1053_),
    .A2(_1079_),
    .B(_1080_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5759_ (.I(_1034_),
    .Z(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5760_ (.I(\as2650.pc[3] ),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5761_ (.I(_1082_),
    .Z(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5762_ (.I(_1083_),
    .Z(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5763_ (.A1(_1084_),
    .A2(_1059_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5764_ (.A1(_0598_),
    .A2(_1081_),
    .B(_1085_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5765_ (.I(_1086_),
    .Z(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5766_ (.A1(\as2650.stack[1][3] ),
    .A2(_1063_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5767_ (.A1(_1053_),
    .A2(_1087_),
    .B(_1088_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5768_ (.I(_1052_),
    .Z(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5769_ (.I(_0699_),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5770_ (.I(\as2650.pc[4] ),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5771_ (.I0(_1090_),
    .I1(_1091_),
    .S(_1009_),
    .Z(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5772_ (.I(_1092_),
    .Z(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5773_ (.I(_1052_),
    .Z(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5774_ (.A1(\as2650.stack[1][4] ),
    .A2(_1094_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5775_ (.A1(_1089_),
    .A2(_1093_),
    .B(_1095_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5776_ (.I(\as2650.pc[5] ),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5777_ (.I(_1096_),
    .Z(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5778_ (.A1(_1097_),
    .A2(_1059_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5779_ (.A1(_0784_),
    .A2(_1081_),
    .B(_1098_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5780_ (.I(_1099_),
    .Z(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5781_ (.A1(\as2650.stack[1][5] ),
    .A2(_1094_),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5782_ (.A1(_1089_),
    .A2(_1100_),
    .B(_1101_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5783_ (.I(_0823_),
    .Z(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5784_ (.I(\as2650.pc[6] ),
    .Z(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5785_ (.I(_1103_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5786_ (.I(_1104_),
    .Z(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5787_ (.A1(_1105_),
    .A2(_0974_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5788_ (.A1(_1102_),
    .A2(_1081_),
    .B(_1106_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5789_ (.I(_1107_),
    .Z(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5790_ (.A1(\as2650.stack[1][6] ),
    .A2(_1094_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5791_ (.A1(_1089_),
    .A2(_1108_),
    .B(_1109_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5792_ (.I(\as2650.pc[7] ),
    .Z(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5793_ (.I(_1110_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5794_ (.I(_1111_),
    .Z(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5795_ (.A1(_1112_),
    .A2(_0974_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5796_ (.A1(_0862_),
    .A2(_1081_),
    .B(_1113_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5797_ (.I(_1114_),
    .Z(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5798_ (.A1(\as2650.stack[1][7] ),
    .A2(_1094_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5799_ (.A1(_1089_),
    .A2(_1115_),
    .B(_1116_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5800_ (.I(_0955_),
    .Z(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5801_ (.I(_1117_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5802_ (.A1(_1046_),
    .A2(_1048_),
    .A3(_1118_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5803_ (.I(_1119_),
    .Z(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5804_ (.I(_1119_),
    .Z(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5805_ (.A1(\as2650.stack[0][0] ),
    .A2(_1121_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5806_ (.A1(_1062_),
    .A2(_1120_),
    .B(_1122_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5807_ (.A1(\as2650.stack[0][1] ),
    .A2(_1121_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5808_ (.A1(_1071_),
    .A2(_1120_),
    .B(_1123_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5809_ (.A1(\as2650.stack[0][2] ),
    .A2(_1121_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5810_ (.A1(_1079_),
    .A2(_1120_),
    .B(_1124_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5811_ (.A1(\as2650.stack[0][3] ),
    .A2(_1121_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5812_ (.A1(_1087_),
    .A2(_1120_),
    .B(_1125_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5813_ (.I(_1119_),
    .Z(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5814_ (.I(_1119_),
    .Z(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5815_ (.A1(\as2650.stack[0][4] ),
    .A2(_1127_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5816_ (.A1(_1093_),
    .A2(_1126_),
    .B(_1128_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5817_ (.A1(\as2650.stack[0][5] ),
    .A2(_1127_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5818_ (.A1(_1100_),
    .A2(_1126_),
    .B(_1129_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5819_ (.A1(\as2650.stack[0][6] ),
    .A2(_1127_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5820_ (.A1(_1108_),
    .A2(_1126_),
    .B(_1130_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5821_ (.A1(\as2650.stack[0][7] ),
    .A2(_1127_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5822_ (.A1(_1115_),
    .A2(_1126_),
    .B(_1131_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5823_ (.I(\as2650.r123_2[3][0] ),
    .Z(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5824_ (.I(_1132_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5825_ (.I(\as2650.r123_2[3][1] ),
    .Z(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5826_ (.I(_1133_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5827_ (.I(\as2650.r123_2[3][2] ),
    .Z(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5828_ (.I(_1134_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5829_ (.I(\as2650.r123_2[3][3] ),
    .Z(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5830_ (.I(_1135_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5831_ (.I(\as2650.r123_2[3][4] ),
    .Z(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5832_ (.I(_1136_),
    .Z(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5833_ (.I(\as2650.r123_2[3][5] ),
    .Z(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5834_ (.I(_1137_),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5835_ (.I(\as2650.r123_2[3][6] ),
    .Z(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5836_ (.I(_1138_),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5837_ (.I(\as2650.r123_2[3][7] ),
    .Z(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5838_ (.I(_1139_),
    .Z(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5839_ (.A1(_0496_),
    .A2(_0919_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5840_ (.A1(_1140_),
    .A2(_1049_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5841_ (.I(_1141_),
    .Z(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5842_ (.I(_1142_),
    .Z(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5843_ (.I(_1142_),
    .Z(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5844_ (.A1(\as2650.stack[1][8] ),
    .A2(_1144_),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5845_ (.A1(_0977_),
    .A2(_1143_),
    .B(_1145_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5846_ (.I(_1141_),
    .Z(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5847_ (.A1(\as2650.stack[1][9] ),
    .A2(_1146_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5848_ (.A1(_0990_),
    .A2(_1143_),
    .B(_1147_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5849_ (.A1(\as2650.stack[1][10] ),
    .A2(_1146_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5850_ (.A1(_1001_),
    .A2(_1143_),
    .B(_1148_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5851_ (.A1(\as2650.stack[1][11] ),
    .A2(_1146_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5852_ (.A1(_1012_),
    .A2(_1143_),
    .B(_1149_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5853_ (.A1(\as2650.stack[1][12] ),
    .A2(_1146_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5854_ (.A1(_1021_),
    .A2(_1144_),
    .B(_1150_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5855_ (.A1(\as2650.stack[1][13] ),
    .A2(_1142_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5856_ (.A1(_1028_),
    .A2(_1144_),
    .B(_1151_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5857_ (.A1(\as2650.stack[1][14] ),
    .A2(_1142_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5858_ (.A1(_1043_),
    .A2(_1144_),
    .B(_1152_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5859_ (.I(\as2650.r123_2[0][0] ),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5860_ (.I(_0332_),
    .Z(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5861_ (.I(_1154_),
    .Z(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5862_ (.A1(_4113_),
    .A2(_4172_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5863_ (.A1(_1155_),
    .A2(_1156_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5864_ (.A1(_4177_),
    .A2(_1156_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5865_ (.A1(_4186_),
    .A2(_4229_),
    .A3(_1158_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5866_ (.I(_1159_),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5867_ (.A1(_4441_),
    .A2(_4412_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5868_ (.A1(_1160_),
    .A2(_1161_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5869_ (.A1(_4220_),
    .A2(_4125_),
    .A3(_1158_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5870_ (.I(_1163_),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5871_ (.I(_1164_),
    .Z(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5872_ (.I(_4263_),
    .Z(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5873_ (.A1(_4233_),
    .A2(_4227_),
    .A3(_4372_),
    .A4(_4277_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5874_ (.A1(_0935_),
    .A2(_1166_),
    .A3(_1167_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5875_ (.A1(_4403_),
    .A2(_4117_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5876_ (.I(_1169_),
    .Z(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5877_ (.A1(_1168_),
    .A2(_1170_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5878_ (.A1(_4166_),
    .A2(_1169_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5879_ (.A1(_4250_),
    .A2(_1172_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5880_ (.A1(_4247_),
    .A2(_1173_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5881_ (.A1(_4268_),
    .A2(_4446_),
    .A3(_1173_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5882_ (.A1(_1165_),
    .A2(_1171_),
    .A3(_1174_),
    .A4(_1175_),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _5883_ (.A1(_4204_),
    .A2(_1158_),
    .B(_1162_),
    .C(_1176_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5884_ (.A1(_4171_),
    .A2(_1177_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5885_ (.A1(_4170_),
    .A2(_1157_),
    .B(_1178_),
    .C(_4284_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5886_ (.I(_1179_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5887_ (.I(_1180_),
    .Z(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5888_ (.A1(_4170_),
    .A2(_1157_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5889_ (.A1(_0332_),
    .A2(_0696_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5890_ (.A1(_1170_),
    .A2(_1183_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5891_ (.A1(_1182_),
    .A2(_1184_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5892_ (.I(_1185_),
    .Z(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5893_ (.I(_4168_),
    .Z(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5894_ (.I(_0945_),
    .Z(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5895_ (.I(_1188_),
    .Z(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5896_ (.A1(_1187_),
    .A2(_1189_),
    .A3(_1156_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5897_ (.I0(_1054_),
    .I1(_4501_),
    .S(_1190_),
    .Z(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5898_ (.I(_1171_),
    .Z(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5899_ (.I(_1175_),
    .Z(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5900_ (.I(_1174_),
    .Z(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5901_ (.I(_1194_),
    .Z(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5902_ (.I(_1160_),
    .Z(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5903_ (.I(_4166_),
    .Z(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5904_ (.A1(_4441_),
    .A2(_1197_),
    .A3(_4221_),
    .A4(_4214_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5905_ (.I(_1198_),
    .Z(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5906_ (.I(_4384_),
    .Z(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5907_ (.I(_1164_),
    .Z(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5908_ (.I(_1198_),
    .Z(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5909_ (.I(net6),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5910_ (.A1(_4394_),
    .A2(_1158_),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5911_ (.I(_1204_),
    .Z(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5912_ (.I(_4216_),
    .Z(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5913_ (.A1(_1206_),
    .A2(_0931_),
    .A3(_4201_),
    .A4(_1172_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5914_ (.I(_1207_),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5915_ (.I(_1163_),
    .Z(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5916_ (.A1(_1203_),
    .A2(_1205_),
    .B1(_1208_),
    .B2(_4399_),
    .C(_1209_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5917_ (.A1(_1200_),
    .A2(_1201_),
    .B(_1202_),
    .C(_1210_),
    .ZN(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5918_ (.I(_1160_),
    .Z(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5919_ (.A1(_4371_),
    .A2(_1199_),
    .B(_1211_),
    .C(_1212_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5920_ (.A1(_4354_),
    .A2(_1196_),
    .B(_1194_),
    .C(_1213_),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5921_ (.A1(_4438_),
    .A2(_1195_),
    .B(_1193_),
    .C(_1214_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5922_ (.A1(_4459_),
    .A2(_1193_),
    .B(_1215_),
    .C(_1192_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5923_ (.A1(_4347_),
    .A2(_1192_),
    .B(_1216_),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5924_ (.I(_1178_),
    .Z(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5925_ (.I(_1218_),
    .Z(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5926_ (.I(_1179_),
    .Z(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5927_ (.A1(_1186_),
    .A2(_1191_),
    .B1(_1217_),
    .B2(_1219_),
    .C(_1220_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5928_ (.A1(_1153_),
    .A2(_1181_),
    .B(_1221_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5929_ (.I(\as2650.r123_2[0][1] ),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5930_ (.I(_1190_),
    .Z(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5931_ (.I(_1190_),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5932_ (.A1(_1065_),
    .A2(_1224_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5933_ (.A1(_0398_),
    .A2(_1223_),
    .B(_1225_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5934_ (.A1(_4265_),
    .A2(_1170_),
    .Z(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5935_ (.I(_1227_),
    .Z(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5936_ (.I(_4441_),
    .Z(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5937_ (.I(_1197_),
    .Z(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5938_ (.A1(_1229_),
    .A2(_1230_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5939_ (.A1(_4445_),
    .A2(_4448_),
    .A3(_1231_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5940_ (.I(_1159_),
    .Z(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5941_ (.I(_1233_),
    .Z(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5942_ (.I(_1202_),
    .Z(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5943_ (.I(_0350_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5944_ (.I(_1204_),
    .Z(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5945_ (.I(_1237_),
    .Z(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5946_ (.A1(_1236_),
    .A2(_1238_),
    .B1(_1208_),
    .B2(_0361_),
    .C(_1165_),
    .ZN(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5947_ (.A1(_0459_),
    .A2(_1201_),
    .B(_1202_),
    .C(_1239_),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5948_ (.A1(_0368_),
    .A2(_1235_),
    .B(_1240_),
    .C(_1212_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5949_ (.A1(_0330_),
    .A2(_1234_),
    .B(_1194_),
    .C(_1241_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5950_ (.A1(_4248_),
    .A2(_1173_),
    .Z(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5951_ (.A1(_0328_),
    .A2(_1243_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5952_ (.A1(_1242_),
    .A2(_1244_),
    .B(_1232_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5953_ (.A1(_0320_),
    .A2(_1232_),
    .B(_1245_),
    .C(_1227_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5954_ (.A1(_0313_),
    .A2(_1228_),
    .B(_1246_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5955_ (.A1(_1186_),
    .A2(_1226_),
    .B1(_1247_),
    .B2(_1219_),
    .C(_1220_),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5956_ (.A1(_1222_),
    .A2(_1181_),
    .B(_1248_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5957_ (.I(\as2650.r123_2[0][2] ),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5958_ (.A1(_0506_),
    .A2(_1224_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5959_ (.A1(_0505_),
    .A2(_1223_),
    .B(_1250_),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5960_ (.I(_4268_),
    .Z(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _5961_ (.A1(_1229_),
    .A2(_1230_),
    .A3(_1252_),
    .A4(_4279_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5962_ (.I(_0438_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5963_ (.I(_1164_),
    .Z(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5964_ (.A1(_0463_),
    .A2(_1237_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5965_ (.A1(_0456_),
    .A2(_1205_),
    .B(_1256_),
    .C(_1165_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5966_ (.A1(_0452_),
    .A2(_1255_),
    .B(_1202_),
    .C(_1257_),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5967_ (.A1(_1200_),
    .A2(_1199_),
    .B(_1258_),
    .C(_1233_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5968_ (.A1(_1254_),
    .A2(_1196_),
    .B(_1259_),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5969_ (.I0(_0476_),
    .I1(_1260_),
    .S(_1195_),
    .Z(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5970_ (.A1(_4265_),
    .A2(_1170_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5971_ (.A1(_0485_),
    .A2(_1253_),
    .B(_1262_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5972_ (.A1(_1253_),
    .A2(_1261_),
    .B(_1263_),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5973_ (.A1(_0437_),
    .A2(_1228_),
    .B(_1264_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5974_ (.A1(_1186_),
    .A2(_1251_),
    .B1(_1265_),
    .B2(_1218_),
    .C(_1220_),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5975_ (.A1(_1249_),
    .A2(_1181_),
    .B(_1266_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5976_ (.I(\as2650.r123_2[0][3] ),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5977_ (.A1(_0598_),
    .A2(_1224_),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5978_ (.A1(_0597_),
    .A2(_1223_),
    .B(_1268_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5979_ (.A1(_0480_),
    .A2(_0572_),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _5980_ (.A1(_4457_),
    .A2(_0451_),
    .B1(_0570_),
    .B2(_0578_),
    .C(_1270_),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5981_ (.I(_1198_),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5982_ (.A1(_0560_),
    .A2(_1237_),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5983_ (.A1(_0556_),
    .A2(_1205_),
    .B(_1273_),
    .C(_1209_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5984_ (.A1(_0553_),
    .A2(_1255_),
    .B(_1274_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5985_ (.A1(_1272_),
    .A2(_1275_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5986_ (.A1(_0348_),
    .A2(_1235_),
    .B(_1276_),
    .C(_1212_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5987_ (.A1(_0543_),
    .A2(_1234_),
    .B(_1195_),
    .C(_1277_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5988_ (.I(_1243_),
    .Z(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5989_ (.A1(_0575_),
    .A2(_1279_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5990_ (.A1(_1193_),
    .A2(_1278_),
    .A3(_1280_),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5991_ (.A1(_1271_),
    .A2(_1193_),
    .B(_1281_),
    .C(_1192_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5992_ (.A1(_0541_),
    .A2(_1192_),
    .B(_1282_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5993_ (.A1(_1185_),
    .A2(_1269_),
    .B1(_1283_),
    .B2(_1218_),
    .C(_1179_),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5994_ (.A1(_1267_),
    .A2(_1181_),
    .B(_1284_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5995_ (.I(\as2650.r123_2[0][4] ),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5996_ (.I(_1180_),
    .Z(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5997_ (.A1(_4442_),
    .A2(_1230_),
    .A3(_1252_),
    .A4(_4279_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5998_ (.I(_0675_),
    .Z(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5999_ (.A1(_1288_),
    .A2(_1205_),
    .B1(_1208_),
    .B2(_0673_),
    .C(_1209_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6000_ (.A1(_0664_),
    .A2(_1255_),
    .B(_1289_),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6001_ (.A1(_1272_),
    .A2(_1290_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6002_ (.A1(_0452_),
    .A2(_1235_),
    .B(_1291_),
    .C(_1212_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6003_ (.A1(_0699_),
    .A2(_1234_),
    .B(_1195_),
    .C(_1292_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6004_ (.A1(_0686_),
    .A2(_1279_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6005_ (.A1(_1287_),
    .A2(_1293_),
    .A3(_1294_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6006_ (.A1(_0643_),
    .A2(_1253_),
    .B(_1295_),
    .C(_1262_),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6007_ (.A1(_0634_),
    .A2(_1262_),
    .B(_1296_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6008_ (.I(_1184_),
    .Z(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6009_ (.A1(_0709_),
    .A2(_1157_),
    .B1(_1182_),
    .B2(_1298_),
    .C(_0700_),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6010_ (.A1(_1219_),
    .A2(_1297_),
    .B(_1299_),
    .C(_1180_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6011_ (.A1(_1285_),
    .A2(_1286_),
    .B(_1300_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6012_ (.I(\as2650.r123_2[0][5] ),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6013_ (.A1(_4445_),
    .A2(_4448_),
    .A3(_1231_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6014_ (.A1(_0762_),
    .A2(_1238_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6015_ (.A1(_0758_),
    .A2(_1238_),
    .B(_1303_),
    .C(_1255_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6016_ (.A1(_0754_),
    .A2(_1201_),
    .B(_1199_),
    .C(_1304_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6017_ (.A1(_0742_),
    .A2(_1235_),
    .B(_1305_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6018_ (.A1(_0783_),
    .A2(_1196_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6019_ (.A1(_1234_),
    .A2(_1306_),
    .B(_1307_),
    .C(_1279_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6020_ (.A1(_0741_),
    .A2(_1279_),
    .B(_1302_),
    .C(_1308_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6021_ (.A1(_0771_),
    .A2(_1287_),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6022_ (.A1(_0736_),
    .A2(_1227_),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6023_ (.A1(_1228_),
    .A2(_1309_),
    .A3(_1310_),
    .B(_1311_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6024_ (.A1(_4509_),
    .A2(_0781_),
    .A3(_1157_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6025_ (.A1(_0784_),
    .A2(_4510_),
    .B(_1185_),
    .C(_1313_),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6026_ (.I(_1314_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6027_ (.A1(_1219_),
    .A2(_1312_),
    .B(_1315_),
    .C(_1220_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6028_ (.A1(_1301_),
    .A2(_1286_),
    .B(_1316_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6029_ (.I(\as2650.r123_2[0][6] ),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6030_ (.A1(_0823_),
    .A2(_1224_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6031_ (.A1(_0854_),
    .A2(_1223_),
    .B(_1318_),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6032_ (.A1(_0833_),
    .A2(_1238_),
    .B1(_1208_),
    .B2(_0829_),
    .C(_1165_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6033_ (.A1(_0826_),
    .A2(_1201_),
    .B(_1320_),
    .ZN(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6034_ (.A1(_0664_),
    .A2(_1272_),
    .B(_1160_),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6035_ (.A1(_1199_),
    .A2(_1321_),
    .B(_1322_),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6036_ (.I(_4420_),
    .Z(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6037_ (.A1(_1324_),
    .A2(_4429_),
    .A3(_1172_),
    .B1(_1233_),
    .B2(_0822_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6038_ (.A1(_1323_),
    .A2(_1325_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6039_ (.A1(_0841_),
    .A2(_1243_),
    .B(_1302_),
    .C(_1326_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6040_ (.A1(_0821_),
    .A2(_1175_),
    .B(_1171_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6041_ (.A1(_1327_),
    .A2(_1328_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6042_ (.A1(_0814_),
    .A2(_1171_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6043_ (.A1(_1329_),
    .A2(_1330_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6044_ (.I(_1331_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6045_ (.A1(_1185_),
    .A2(_1319_),
    .B1(_1332_),
    .B2(_1218_),
    .C(_1179_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6046_ (.A1(_1317_),
    .A2(_1286_),
    .B(_1333_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6047_ (.I(\as2650.r123_2[0][7] ),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6048_ (.A1(_0863_),
    .A2(_1186_),
    .B(_1180_),
    .ZN(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6049_ (.I(net3),
    .Z(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6050_ (.A1(_1336_),
    .A2(_1237_),
    .B1(_1207_),
    .B2(_0898_),
    .C(_1164_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6051_ (.A1(_0904_),
    .A2(_1209_),
    .B(_1337_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6052_ (.A1(_1198_),
    .A2(_1338_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6053_ (.A1(_0753_),
    .A2(_1272_),
    .B(_1339_),
    .C(_1233_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6054_ (.A1(_0909_),
    .A2(_1196_),
    .B(_1194_),
    .C(_1340_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6055_ (.A1(_0894_),
    .A2(_1243_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6056_ (.A1(_1175_),
    .A2(_1341_),
    .A3(_1342_),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6057_ (.A1(_0891_),
    .A2(_1253_),
    .B(_1343_),
    .ZN(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6058_ (.A1(_1227_),
    .A2(_1344_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6059_ (.A1(_0883_),
    .A2(_1228_),
    .B(_1345_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6060_ (.A1(_4171_),
    .A2(_1177_),
    .A3(_1346_),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6061_ (.A1(_1334_),
    .A2(_1286_),
    .B1(_1335_),
    .B2(_1347_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6062_ (.I(_4158_),
    .Z(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6063_ (.I(_4226_),
    .Z(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6064_ (.I(_0333_),
    .Z(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6065_ (.I(_1350_),
    .Z(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6066_ (.A1(_1349_),
    .A2(_1351_),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6067_ (.I(_4362_),
    .Z(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6068_ (.A1(\as2650.psl[7] ),
    .A2(_4150_),
    .Z(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6069_ (.A1(\as2650.psl[6] ),
    .A2(_4367_),
    .Z(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6070_ (.A1(_1354_),
    .A2(_1355_),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _6071_ (.A1(_4157_),
    .A2(_1353_),
    .A3(_1356_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6072_ (.A1(_1348_),
    .A2(_1357_),
    .B(_0930_),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6073_ (.A1(_0921_),
    .A2(_4291_),
    .A3(_4138_),
    .ZN(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6074_ (.A1(_0921_),
    .A2(_0670_),
    .ZN(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6075_ (.A1(_1359_),
    .A2(_1360_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6076_ (.A1(_4209_),
    .A2(_4157_),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6077_ (.A1(_4200_),
    .A2(_1362_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6078_ (.A1(_1361_),
    .A2(_1363_),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6079_ (.A1(_4405_),
    .A2(_1364_),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6080_ (.A1(_4367_),
    .A2(_4150_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6081_ (.I(_1366_),
    .Z(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6082_ (.I(_4390_),
    .Z(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6083_ (.A1(_0922_),
    .A2(_1368_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6084_ (.A1(_4292_),
    .A2(_4199_),
    .A3(_1369_),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6085_ (.I(_1370_),
    .Z(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6086_ (.I(_0931_),
    .Z(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6087_ (.I(_1372_),
    .Z(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6088_ (.A1(_1367_),
    .A2(_1371_),
    .B(_1364_),
    .C(_1373_),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6089_ (.A1(_4221_),
    .A2(_4514_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6090_ (.I(_0694_),
    .Z(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6091_ (.A1(_4206_),
    .A2(_1376_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6092_ (.I(_4114_),
    .Z(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6093_ (.A1(_1368_),
    .A2(_4181_),
    .ZN(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6094_ (.I(_1379_),
    .Z(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6095_ (.A1(_4210_),
    .A2(_1206_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _6096_ (.A1(_0294_),
    .A2(_4420_),
    .A3(_4218_),
    .A4(_1381_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6097_ (.A1(_0693_),
    .A2(_1382_),
    .ZN(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6098_ (.I(_4191_),
    .Z(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6099_ (.A1(_4192_),
    .A2(_4404_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6100_ (.A1(_1384_),
    .A2(_1385_),
    .ZN(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6101_ (.I(_1386_),
    .Z(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6102_ (.I(_1387_),
    .Z(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6103_ (.A1(_0922_),
    .A2(_4181_),
    .A3(_4294_),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6104_ (.A1(_1388_),
    .A2(_1389_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6105_ (.A1(_1378_),
    .A2(_1380_),
    .A3(_1383_),
    .A4(_1390_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6106_ (.A1(_1375_),
    .A2(_1377_),
    .A3(_1391_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6107_ (.A1(_1365_),
    .A2(_1374_),
    .A3(_1392_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6108_ (.I(_4206_),
    .Z(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6109_ (.I(_1394_),
    .Z(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6110_ (.I(_4219_),
    .Z(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6111_ (.A1(_1396_),
    .A2(_4213_),
    .ZN(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6112_ (.I(_1397_),
    .Z(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6113_ (.A1(_0697_),
    .A2(_1398_),
    .ZN(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6114_ (.I(_4132_),
    .Z(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6115_ (.A1(_4171_),
    .A2(_1400_),
    .A3(_1348_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6116_ (.A1(_0946_),
    .A2(_1401_),
    .Z(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6117_ (.A1(_0691_),
    .A2(_0692_),
    .ZN(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6118_ (.A1(_4133_),
    .A2(_4145_),
    .A3(_1403_),
    .ZN(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6119_ (.A1(_1402_),
    .A2(_1404_),
    .Z(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6120_ (.A1(_1395_),
    .A2(_1363_),
    .A3(_1399_),
    .A4(_1405_),
    .ZN(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6121_ (.A1(_1358_),
    .A2(_1393_),
    .A3(_1406_),
    .ZN(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6122_ (.A1(_4391_),
    .A2(_1361_),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6123_ (.A1(_1348_),
    .A2(_1352_),
    .B(_1407_),
    .C(_1408_),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6124_ (.I(_0758_),
    .Z(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6125_ (.I(_1410_),
    .Z(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6126_ (.A1(_1230_),
    .A2(_1382_),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6127_ (.I(_1412_),
    .Z(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6128_ (.A1(\as2650.psu[5] ),
    .A2(_1411_),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6129_ (.I(_1387_),
    .Z(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6130_ (.I(_1415_),
    .Z(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6131_ (.I(_1416_),
    .Z(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6132_ (.A1(_1411_),
    .A2(_1413_),
    .B(_1414_),
    .C(_1417_),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6133_ (.I(_0333_),
    .Z(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6134_ (.I(_1419_),
    .Z(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6135_ (.A1(_0651_),
    .A2(_1420_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6136_ (.I(_1389_),
    .Z(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6137_ (.A1(_1418_),
    .A2(_1421_),
    .B(_1422_),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6138_ (.I(_4116_),
    .Z(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6139_ (.I(_1424_),
    .Z(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6140_ (.A1(\as2650.psu[5] ),
    .A2(_1409_),
    .B(_1425_),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6141_ (.A1(_1409_),
    .A2(_1423_),
    .B(_1426_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6142_ (.I(_4284_),
    .Z(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6143_ (.I(_1427_),
    .Z(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6144_ (.I(\as2650.psl[6] ),
    .Z(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6145_ (.I(_1365_),
    .ZN(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6146_ (.A1(_0930_),
    .A2(_1388_),
    .A3(_0696_),
    .A4(_1389_),
    .ZN(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6147_ (.A1(_1430_),
    .A2(_1431_),
    .B(_1380_),
    .ZN(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6148_ (.A1(_1368_),
    .A2(_1397_),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6149_ (.A1(_4186_),
    .A2(_1433_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6150_ (.I(_4143_),
    .Z(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6151_ (.A1(_1435_),
    .A2(_4200_),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6152_ (.A1(_4185_),
    .A2(_1436_),
    .ZN(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6153_ (.A1(_1183_),
    .A2(_1434_),
    .A3(_1437_),
    .ZN(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6154_ (.A1(_4311_),
    .A2(_4410_),
    .A3(_1374_),
    .ZN(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6155_ (.A1(_1438_),
    .A2(_1439_),
    .ZN(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6156_ (.A1(_4232_),
    .A2(_4167_),
    .A3(_4340_),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6157_ (.I(_4193_),
    .Z(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6158_ (.I(_4124_),
    .Z(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6159_ (.A1(_4393_),
    .A2(_1441_),
    .B(_1442_),
    .C(_1443_),
    .ZN(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6160_ (.A1(_4233_),
    .A2(_4126_),
    .ZN(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6161_ (.I(_1445_),
    .Z(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6162_ (.A1(_4372_),
    .A2(_4406_),
    .A3(_0335_),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6163_ (.A1(_4124_),
    .A2(_4202_),
    .B(_1447_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6164_ (.A1(_1400_),
    .A2(_1446_),
    .B(_1448_),
    .ZN(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6165_ (.I(_4233_),
    .Z(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6166_ (.A1(_1450_),
    .A2(_0945_),
    .ZN(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6167_ (.A1(_0935_),
    .A2(_1372_),
    .ZN(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6168_ (.A1(_1451_),
    .A2(_1452_),
    .ZN(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6169_ (.I(_0691_),
    .Z(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6170_ (.I(_0931_),
    .Z(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6171_ (.I(_1455_),
    .Z(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6172_ (.A1(_1454_),
    .A2(_1456_),
    .A3(_1382_),
    .ZN(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6173_ (.I(_4225_),
    .Z(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6174_ (.I(_4123_),
    .Z(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6175_ (.I(_4252_),
    .Z(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6176_ (.A1(_1459_),
    .A2(_1460_),
    .ZN(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6177_ (.A1(_1458_),
    .A2(_1372_),
    .B(_1461_),
    .ZN(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6178_ (.I(_1462_),
    .Z(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6179_ (.A1(_1449_),
    .A2(_1453_),
    .A3(_1457_),
    .A4(_1463_),
    .ZN(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6180_ (.I(_4222_),
    .Z(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6181_ (.I(_1465_),
    .Z(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6182_ (.A1(_1349_),
    .A2(_4513_),
    .A3(_0655_),
    .ZN(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6183_ (.I(_4294_),
    .Z(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6184_ (.A1(_4154_),
    .A2(_4225_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6185_ (.A1(_1468_),
    .A2(_1469_),
    .ZN(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6186_ (.A1(_1441_),
    .A2(_1470_),
    .ZN(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6187_ (.A1(_1445_),
    .A2(_1471_),
    .ZN(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6188_ (.A1(_1384_),
    .A2(_4237_),
    .ZN(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6189_ (.A1(_4114_),
    .A2(_1473_),
    .ZN(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6190_ (.I(_1368_),
    .Z(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6191_ (.I(_1450_),
    .Z(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6192_ (.A1(_1475_),
    .A2(_1476_),
    .ZN(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6193_ (.A1(_4465_),
    .A2(_0971_),
    .B(_1154_),
    .ZN(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6194_ (.A1(_1477_),
    .A2(_1478_),
    .ZN(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6195_ (.A1(_1422_),
    .A2(_1377_),
    .A3(_1474_),
    .A4(_1479_),
    .ZN(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6196_ (.A1(_1466_),
    .A2(_1467_),
    .B1(_1472_),
    .B2(_0335_),
    .C(_1480_),
    .ZN(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6197_ (.A1(_1464_),
    .A2(_1481_),
    .ZN(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6198_ (.A1(_1432_),
    .A2(_1440_),
    .A3(_1444_),
    .A4(_1482_),
    .ZN(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6199_ (.A1(_1429_),
    .A2(_1483_),
    .ZN(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6200_ (.A1(_1458_),
    .A2(_1387_),
    .ZN(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6201_ (.I(_1485_),
    .Z(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6202_ (.I(_1486_),
    .Z(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6203_ (.I(_1487_),
    .Z(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6204_ (.A1(_4347_),
    .A2(_0541_),
    .A3(_0633_),
    .ZN(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6205_ (.A1(_0313_),
    .A2(_0437_),
    .A3(_0814_),
    .ZN(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6206_ (.A1(_0736_),
    .A2(_1489_),
    .A3(_1490_),
    .ZN(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6207_ (.I(\as2650.psl[1] ),
    .Z(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6208_ (.I(_0873_),
    .Z(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6209_ (.I(_0870_),
    .ZN(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6210_ (.A1(_0721_),
    .A2(_0723_),
    .B(_0806_),
    .ZN(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6211_ (.A1(_0799_),
    .A2(_0797_),
    .ZN(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6212_ (.A1(_0802_),
    .A2(_1495_),
    .B(_1496_),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6213_ (.A1(_1493_),
    .A2(_1497_),
    .ZN(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6214_ (.A1(_0866_),
    .A2(_1494_),
    .B(_1498_),
    .ZN(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6215_ (.A1(_0301_),
    .A2(_0290_),
    .ZN(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6216_ (.A1(_0432_),
    .A2(_0419_),
    .B1(_0423_),
    .B2(_1500_),
    .ZN(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6217_ (.A1(_0526_),
    .A2(_1501_),
    .B(_0532_),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6218_ (.A1(_0621_),
    .A2(_0722_),
    .A3(_0801_),
    .A4(_1493_),
    .ZN(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6219_ (.A1(_0623_),
    .A2(_1502_),
    .B(_1503_),
    .ZN(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6220_ (.A1(_1492_),
    .A2(_1493_),
    .B1(_1499_),
    .B2(_1504_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6221_ (.A1(_1492_),
    .A2(_1493_),
    .A3(_1499_),
    .B(_1505_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6222_ (.A1(_1166_),
    .A2(_1506_),
    .ZN(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6223_ (.A1(_4330_),
    .A2(_0291_),
    .A3(_0421_),
    .A4(_0532_),
    .ZN(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6224_ (.A1(_1503_),
    .A2(_1508_),
    .ZN(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6225_ (.A1(_1166_),
    .A2(_0884_),
    .A3(_1491_),
    .B1(_1507_),
    .B2(_1509_),
    .ZN(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6226_ (.I(_1458_),
    .Z(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6227_ (.I(_1511_),
    .Z(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6228_ (.I(_1512_),
    .Z(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6229_ (.I(_4201_),
    .Z(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6230_ (.I(_1514_),
    .Z(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6231_ (.A1(_1360_),
    .A2(_4371_),
    .ZN(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6232_ (.I(_1360_),
    .Z(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6233_ (.A1(_1517_),
    .A2(_0792_),
    .ZN(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6234_ (.I(_4213_),
    .Z(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6235_ (.I(_1519_),
    .Z(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6236_ (.I(_1369_),
    .Z(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6237_ (.I(_1521_),
    .Z(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6238_ (.I(_4251_),
    .Z(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6239_ (.A1(_1523_),
    .A2(_0969_),
    .ZN(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6240_ (.I(_0832_),
    .Z(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6241_ (.A1(_0692_),
    .A2(_0833_),
    .ZN(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6242_ (.A1(_1429_),
    .A2(_1525_),
    .B(_0431_),
    .C(_1526_),
    .ZN(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6243_ (.A1(_4148_),
    .A2(_1522_),
    .A3(_1524_),
    .A4(_1527_),
    .ZN(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6244_ (.A1(_0438_),
    .A2(_0330_),
    .A3(_4353_),
    .ZN(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6245_ (.A1(_0822_),
    .A2(_0783_),
    .A3(_0644_),
    .A4(_0519_),
    .ZN(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6246_ (.A1(_1529_),
    .A2(_1530_),
    .B(_0860_),
    .ZN(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6247_ (.A1(_1401_),
    .A2(_1531_),
    .ZN(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6248_ (.A1(_0793_),
    .A2(_1401_),
    .B(_1532_),
    .C(_1419_),
    .ZN(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6249_ (.A1(_1528_),
    .A2(_1533_),
    .ZN(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6250_ (.I(_1359_),
    .Z(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6251_ (.A1(_1520_),
    .A2(_1534_),
    .B(_1535_),
    .ZN(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6252_ (.A1(_0815_),
    .A2(_1516_),
    .B(_1518_),
    .C(_1536_),
    .ZN(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6253_ (.I(_1535_),
    .Z(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6254_ (.I(_0754_),
    .Z(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6255_ (.A1(_0827_),
    .A2(_0640_),
    .A3(_0665_),
    .A4(_1539_),
    .ZN(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6256_ (.A1(_1538_),
    .A2(_0905_),
    .A3(_1540_),
    .ZN(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6257_ (.A1(_1515_),
    .A2(_1537_),
    .A3(_1541_),
    .ZN(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6258_ (.I(_1336_),
    .Z(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6259_ (.I(_1543_),
    .Z(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6260_ (.I(_1544_),
    .Z(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6261_ (.I(_4392_),
    .Z(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6262_ (.A1(_1545_),
    .A2(_1546_),
    .ZN(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6263_ (.I(_4392_),
    .Z(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6264_ (.I(_4387_),
    .Z(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6265_ (.I(_1549_),
    .Z(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6266_ (.I(_0353_),
    .Z(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6267_ (.I(_0456_),
    .Z(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6268_ (.I(_1552_),
    .Z(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6269_ (.I(_0555_),
    .Z(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6270_ (.I(_1554_),
    .Z(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6271_ (.I(_1555_),
    .Z(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6272_ (.A1(_1550_),
    .A2(_1551_),
    .A3(_1553_),
    .A4(_1556_),
    .ZN(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6273_ (.I(_0677_),
    .Z(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6274_ (.I(_1525_),
    .Z(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6275_ (.I(_1559_),
    .Z(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6276_ (.A1(_1558_),
    .A2(_1410_),
    .A3(_1560_),
    .ZN(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6277_ (.A1(_1548_),
    .A2(_1557_),
    .A3(_1561_),
    .ZN(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6278_ (.A1(_1513_),
    .A2(_1542_),
    .A3(_1547_),
    .A4(_1562_),
    .ZN(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6279_ (.A1(_1324_),
    .A2(_1419_),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6280_ (.A1(_1468_),
    .A2(_1469_),
    .Z(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6281_ (.A1(_0827_),
    .A2(_0887_),
    .A3(_1565_),
    .ZN(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6282_ (.A1(_1531_),
    .A2(_1470_),
    .ZN(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6283_ (.A1(_1566_),
    .A2(_1567_),
    .ZN(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6284_ (.A1(_1564_),
    .A2(_1568_),
    .ZN(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6285_ (.A1(_1563_),
    .A2(_1569_),
    .A3(_1483_),
    .ZN(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6286_ (.A1(_1488_),
    .A2(_1510_),
    .B(_1570_),
    .ZN(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6287_ (.A1(_1428_),
    .A2(_1484_),
    .A3(_1571_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6288_ (.I(_1512_),
    .Z(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6289_ (.I(_1572_),
    .Z(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6290_ (.I(_1514_),
    .Z(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6291_ (.I(_1396_),
    .Z(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6292_ (.I(_1361_),
    .Z(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6293_ (.I(_1394_),
    .Z(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6294_ (.A1(_4151_),
    .A2(_1370_),
    .ZN(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6295_ (.A1(_1458_),
    .A2(_4333_),
    .ZN(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6296_ (.A1(_1454_),
    .A2(_1579_),
    .A3(_1521_),
    .ZN(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6297_ (.I(_0933_),
    .Z(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6298_ (.I(_0378_),
    .Z(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6299_ (.I(net27),
    .ZN(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6300_ (.I(_0755_),
    .ZN(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6301_ (.I(_1584_),
    .Z(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6302_ (.A1(_4477_),
    .A2(_1236_),
    .B1(_1585_),
    .B2(\as2650.psu[5] ),
    .ZN(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6303_ (.A1(_1582_),
    .A2(_4387_),
    .B1(_0832_),
    .B2(_1583_),
    .C(_1586_),
    .ZN(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6304_ (.I(\as2650.psu[3] ),
    .ZN(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6305_ (.I(\as2650.psu[4] ),
    .ZN(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6306_ (.I(_4486_),
    .Z(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6307_ (.A1(_1588_),
    .A2(_1554_),
    .B1(_0676_),
    .B2(_1589_),
    .C1(_1590_),
    .C2(_0455_),
    .ZN(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6308_ (.A1(\as2650.psu[7] ),
    .A2(_1581_),
    .B(_1587_),
    .C(_1591_),
    .ZN(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6309_ (.A1(_0455_),
    .A2(_0347_),
    .B1(_0451_),
    .B2(_1554_),
    .ZN(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6310_ (.A1(_0691_),
    .A2(_4182_),
    .A3(_4332_),
    .A4(_1381_),
    .ZN(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6311_ (.I(net2),
    .Z(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6312_ (.I(_1595_),
    .Z(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6313_ (.I(_1596_),
    .Z(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6314_ (.A1(_0676_),
    .A2(_0553_),
    .B1(_0664_),
    .B2(_0757_),
    .C1(_0753_),
    .C2(_1597_),
    .ZN(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6315_ (.I(net3),
    .Z(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6316_ (.A1(_4387_),
    .A2(_0367_),
    .B1(_0441_),
    .B2(_0351_),
    .C1(_0826_),
    .C2(_1599_),
    .ZN(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6317_ (.A1(_1593_),
    .A2(_1594_),
    .A3(_1598_),
    .A4(_1600_),
    .Z(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6318_ (.I(\as2650.psl[5] ),
    .ZN(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6319_ (.A1(_4335_),
    .A2(_4386_),
    .B1(_0757_),
    .B2(_1602_),
    .ZN(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6320_ (.I(\as2650.psl[1] ),
    .ZN(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6321_ (.I(_1429_),
    .ZN(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6322_ (.A1(_1604_),
    .A2(_0350_),
    .B1(_1597_),
    .B2(_1605_),
    .ZN(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6323_ (.I(\as2650.psl[3] ),
    .ZN(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6324_ (.I(\as2650.psl[7] ),
    .Z(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6325_ (.I(_0454_),
    .ZN(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6326_ (.A1(_1608_),
    .A2(_0933_),
    .B1(_1609_),
    .B2(\as2650.overflow ),
    .ZN(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6327_ (.A1(_1607_),
    .A2(_0555_),
    .B1(_0675_),
    .B2(_4403_),
    .C(_1610_),
    .ZN(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6328_ (.A1(_1603_),
    .A2(_1606_),
    .A3(_1611_),
    .ZN(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6329_ (.A1(_1454_),
    .A2(_1612_),
    .B(_1521_),
    .C(_1579_),
    .ZN(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6330_ (.A1(_1601_),
    .A2(_1613_),
    .ZN(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6331_ (.A1(_1353_),
    .A2(_1371_),
    .B1(_1580_),
    .B2(_1592_),
    .C(_1614_),
    .ZN(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6332_ (.I(_0901_),
    .Z(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6333_ (.A1(_1608_),
    .A2(_1616_),
    .A3(_1367_),
    .A4(_1382_),
    .ZN(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6334_ (.A1(_1615_),
    .A2(_1617_),
    .ZN(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6335_ (.I(_1608_),
    .ZN(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6336_ (.I(_1336_),
    .Z(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6337_ (.I(_1620_),
    .Z(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6338_ (.A1(_1619_),
    .A2(_1621_),
    .A3(_1578_),
    .ZN(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6339_ (.A1(_1578_),
    .A2(_1618_),
    .B(_1622_),
    .ZN(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6340_ (.I(_1388_),
    .Z(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6341_ (.A1(_0861_),
    .A2(_1624_),
    .ZN(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6342_ (.A1(_1577_),
    .A2(_1623_),
    .B(_1625_),
    .ZN(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6343_ (.A1(_1576_),
    .A2(_1626_),
    .ZN(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6344_ (.A1(_1575_),
    .A2(_0905_),
    .B(_1518_),
    .C(_1627_),
    .ZN(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6345_ (.A1(_1574_),
    .A2(_1628_),
    .ZN(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6346_ (.A1(_1573_),
    .A2(_1547_),
    .A3(_1629_),
    .ZN(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6347_ (.I(_1476_),
    .Z(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6348_ (.I(_1631_),
    .Z(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6349_ (.I(_0970_),
    .Z(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6350_ (.I(_1633_),
    .Z(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6351_ (.A1(_1166_),
    .A2(_0883_),
    .B(_1507_),
    .C(_1634_),
    .ZN(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6352_ (.I(_0827_),
    .Z(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6353_ (.A1(_1636_),
    .A2(_1565_),
    .ZN(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6354_ (.I(_1415_),
    .Z(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6355_ (.I(_1638_),
    .Z(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6356_ (.A1(_0861_),
    .A2(_1565_),
    .B(_1637_),
    .C(_1639_),
    .ZN(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6357_ (.A1(_1632_),
    .A2(_1635_),
    .A3(_1640_),
    .ZN(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6358_ (.A1(_1630_),
    .A2(_1641_),
    .ZN(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6359_ (.A1(_1608_),
    .A2(_1483_),
    .ZN(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6360_ (.I(_1427_),
    .Z(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6361_ (.A1(_1483_),
    .A2(_1642_),
    .B(_1643_),
    .C(_1644_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6362_ (.A1(_1045_),
    .A2(_1047_),
    .A3(_1117_),
    .ZN(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6363_ (.I(_1645_),
    .Z(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6364_ (.I(_1646_),
    .Z(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6365_ (.I(_1646_),
    .Z(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6366_ (.A1(\as2650.stack[6][8] ),
    .A2(_1648_),
    .ZN(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6367_ (.A1(_0977_),
    .A2(_1647_),
    .B(_1649_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6368_ (.I(_1645_),
    .Z(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6369_ (.A1(\as2650.stack[6][9] ),
    .A2(_1650_),
    .ZN(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6370_ (.A1(_0990_),
    .A2(_1647_),
    .B(_1651_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6371_ (.A1(\as2650.stack[6][10] ),
    .A2(_1650_),
    .ZN(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6372_ (.A1(_1001_),
    .A2(_1647_),
    .B(_1652_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6373_ (.A1(\as2650.stack[6][11] ),
    .A2(_1650_),
    .ZN(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6374_ (.A1(_1012_),
    .A2(_1647_),
    .B(_1653_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6375_ (.A1(\as2650.stack[6][12] ),
    .A2(_1650_),
    .ZN(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6376_ (.A1(_1021_),
    .A2(_1648_),
    .B(_1654_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6377_ (.A1(\as2650.stack[6][13] ),
    .A2(_1646_),
    .ZN(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6378_ (.A1(_1028_),
    .A2(_1648_),
    .B(_1655_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6379_ (.A1(\as2650.stack[6][14] ),
    .A2(_1646_),
    .ZN(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6380_ (.A1(_1043_),
    .A2(_1648_),
    .B(_1656_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6381_ (.A1(_1621_),
    .A2(_1456_),
    .ZN(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6382_ (.I(_4405_),
    .Z(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6383_ (.I(_1658_),
    .Z(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6384_ (.A1(_4511_),
    .A2(_1366_),
    .ZN(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6385_ (.A1(_4216_),
    .A2(_1660_),
    .ZN(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6386_ (.A1(_0922_),
    .A2(_1661_),
    .ZN(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6387_ (.I(_1662_),
    .Z(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6388_ (.I(_1663_),
    .Z(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6389_ (.A1(_1659_),
    .A2(_1664_),
    .B(_1473_),
    .ZN(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _6390_ (.A1(_4270_),
    .A2(_1416_),
    .A3(_1657_),
    .A4(_1665_),
    .Z(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6391_ (.I(_1666_),
    .ZN(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6392_ (.I(_1667_),
    .Z(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6393_ (.I(_1550_),
    .Z(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6394_ (.A1(_0943_),
    .A2(_1384_),
    .ZN(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6395_ (.A1(_1442_),
    .A2(_1670_),
    .ZN(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6396_ (.I(_1671_),
    .Z(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6397_ (.I(_1667_),
    .Z(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6398_ (.A1(_4184_),
    .A2(_4225_),
    .ZN(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6399_ (.I(_1674_),
    .Z(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6400_ (.I(_1675_),
    .Z(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6401_ (.I(_1676_),
    .Z(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6402_ (.A1(_1671_),
    .A2(_1677_),
    .ZN(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6403_ (.A1(_1669_),
    .A2(_1672_),
    .B(_1673_),
    .C(_1678_),
    .ZN(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6404_ (.A1(_4148_),
    .A2(_1668_),
    .B(_1679_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6405_ (.I(_0353_),
    .Z(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6406_ (.A1(_1680_),
    .A2(_1672_),
    .B(_1673_),
    .C(_1678_),
    .ZN(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6407_ (.A1(_0692_),
    .A2(_1668_),
    .B(_1681_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6408_ (.I(_0938_),
    .Z(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6409_ (.I(_1553_),
    .Z(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6410_ (.A1(_1672_),
    .A2(_1666_),
    .ZN(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6411_ (.A1(_1683_),
    .A2(_1684_),
    .ZN(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6412_ (.A1(_1682_),
    .A2(_1668_),
    .B(_1685_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6413_ (.A1(_0963_),
    .A2(_1473_),
    .ZN(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6414_ (.I(_1686_),
    .Z(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6415_ (.A1(_1411_),
    .A2(_1672_),
    .B(_1678_),
    .ZN(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6416_ (.A1(_4311_),
    .A2(_1687_),
    .B1(_1688_),
    .B2(_1668_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6417_ (.I(_1560_),
    .Z(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6418_ (.A1(_1689_),
    .A2(_1684_),
    .ZN(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6419_ (.A1(_4141_),
    .A2(_1673_),
    .B(_1690_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6420_ (.I(_1545_),
    .Z(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6421_ (.A1(_1691_),
    .A2(_1684_),
    .ZN(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6422_ (.A1(_4196_),
    .A2(_1673_),
    .B(_1692_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6423_ (.I(_4284_),
    .Z(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6424_ (.A1(_1156_),
    .A2(_1375_),
    .ZN(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6425_ (.I(_1454_),
    .Z(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6426_ (.A1(_1695_),
    .A2(_1177_),
    .Z(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6427_ (.I(_1696_),
    .ZN(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6428_ (.A1(_1693_),
    .A2(_1694_),
    .A3(_1697_),
    .ZN(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6429_ (.I(_1698_),
    .Z(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6430_ (.A1(\as2650.r0[0] ),
    .A2(_0960_),
    .Z(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6431_ (.I(_1700_),
    .Z(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6432_ (.I(_1694_),
    .Z(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6433_ (.I(_1702_),
    .Z(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6434_ (.A1(\as2650.r123_2[1][0] ),
    .A2(_1699_),
    .B1(_1701_),
    .B2(_1703_),
    .ZN(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6435_ (.I(_1697_),
    .Z(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6436_ (.A1(_1217_),
    .A2(_1705_),
    .ZN(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6437_ (.A1(_1704_),
    .A2(_1706_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6438_ (.A1(_0329_),
    .A2(_0984_),
    .A3(_1701_),
    .ZN(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6439_ (.A1(_0331_),
    .A2(_0962_),
    .ZN(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6440_ (.A1(_4503_),
    .A2(_0984_),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6441_ (.A1(_1708_),
    .A2(_1709_),
    .ZN(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6442_ (.A1(_1707_),
    .A2(_1710_),
    .Z(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6443_ (.A1(\as2650.r123_2[1][1] ),
    .A2(_1699_),
    .B1(_1711_),
    .B2(_1703_),
    .ZN(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6444_ (.A1(_1247_),
    .A2(_1705_),
    .ZN(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6445_ (.A1(_1712_),
    .A2(_1713_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6446_ (.A1(_0414_),
    .A2(_0962_),
    .ZN(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6447_ (.A1(_4379_),
    .A2(_4316_),
    .A3(_0982_),
    .A4(_0995_),
    .ZN(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6448_ (.A1(_0286_),
    .A2(_0983_),
    .ZN(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6449_ (.I(_0994_),
    .Z(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6450_ (.A1(_4299_),
    .A2(_1717_),
    .ZN(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6451_ (.A1(_1716_),
    .A2(_1718_),
    .ZN(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6452_ (.A1(_1715_),
    .A2(_1719_),
    .ZN(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6453_ (.A1(_1714_),
    .A2(_1720_),
    .ZN(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6454_ (.A1(_1707_),
    .A2(_1721_),
    .Z(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6455_ (.I(_1702_),
    .Z(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6456_ (.A1(\as2650.r123_2[1][2] ),
    .A2(_1699_),
    .B1(_1722_),
    .B2(_1723_),
    .ZN(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6457_ (.A1(_1265_),
    .A2(_1705_),
    .ZN(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6458_ (.A1(_1724_),
    .A2(_1725_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6459_ (.I(_1698_),
    .Z(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6460_ (.A1(_1707_),
    .A2(_1721_),
    .Z(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6461_ (.A1(_4317_),
    .A2(_1005_),
    .ZN(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6462_ (.A1(_0414_),
    .A2(_0961_),
    .A3(_1715_),
    .A4(_1719_),
    .ZN(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6463_ (.A1(_0444_),
    .A2(_0961_),
    .Z(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6464_ (.A1(_0286_),
    .A2(_4316_),
    .A3(_0982_),
    .A4(_0996_),
    .Z(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6465_ (.A1(_0343_),
    .A2(_0286_),
    .A3(_0983_),
    .A4(_0996_),
    .ZN(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6466_ (.A1(_1731_),
    .A2(_1732_),
    .ZN(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6467_ (.I(\as2650.r0[1] ),
    .Z(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6468_ (.A1(_0342_),
    .A2(_1734_),
    .A3(_0982_),
    .A4(_0995_),
    .Z(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6469_ (.A1(_0343_),
    .A2(_0983_),
    .ZN(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6470_ (.A1(_1734_),
    .A2(_1717_),
    .ZN(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6471_ (.A1(_1715_),
    .A2(_1735_),
    .B1(_1736_),
    .B2(_1737_),
    .ZN(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6472_ (.A1(_1733_),
    .A2(_1738_),
    .Z(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6473_ (.A1(_1729_),
    .A2(_1730_),
    .A3(_1739_),
    .Z(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6474_ (.A1(_1728_),
    .A2(_1740_),
    .ZN(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6475_ (.A1(_1727_),
    .A2(_1741_),
    .ZN(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6476_ (.I(_1742_),
    .ZN(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6477_ (.A1(\as2650.r123_2[1][3] ),
    .A2(_1726_),
    .B1(_1743_),
    .B2(_1723_),
    .ZN(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6478_ (.A1(_1283_),
    .A2(_1705_),
    .ZN(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6479_ (.A1(_1744_),
    .A2(_1745_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6480_ (.A1(_1727_),
    .A2(_1741_),
    .ZN(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6481_ (.A1(_1730_),
    .A2(_1739_),
    .ZN(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6482_ (.A1(_1714_),
    .A2(_1720_),
    .A3(_1747_),
    .B1(_1740_),
    .B2(_1728_),
    .ZN(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6483_ (.A1(_0329_),
    .A2(_1004_),
    .ZN(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6484_ (.A1(_1731_),
    .A2(_1732_),
    .B1(_1738_),
    .B2(_1730_),
    .ZN(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6485_ (.A1(_0545_),
    .A2(_0960_),
    .ZN(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6486_ (.I(_0994_),
    .Z(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6487_ (.A1(\as2650.r0[2] ),
    .A2(_1752_),
    .ZN(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6488_ (.A1(_0442_),
    .A2(_0981_),
    .ZN(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6489_ (.A1(_4299_),
    .A2(_1016_),
    .ZN(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6490_ (.A1(_1753_),
    .A2(_1754_),
    .A3(_1755_),
    .ZN(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6491_ (.A1(_1735_),
    .A2(_1751_),
    .A3(_1756_),
    .Z(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6492_ (.A1(_1750_),
    .A2(_1757_),
    .ZN(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6493_ (.A1(_1749_),
    .A2(_1758_),
    .Z(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6494_ (.A1(_1748_),
    .A2(_1759_),
    .Z(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6495_ (.A1(_1746_),
    .A2(_1760_),
    .ZN(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6496_ (.A1(_1298_),
    .A2(_1761_),
    .ZN(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6497_ (.A1(\as2650.r123_2[1][4] ),
    .A2(_1699_),
    .B(_1762_),
    .ZN(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6498_ (.A1(_1297_),
    .A2(_1697_),
    .ZN(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6499_ (.A1(_1763_),
    .A2(_1764_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6500_ (.A1(_1748_),
    .A2(_1759_),
    .Z(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6501_ (.A1(_1746_),
    .A2(_1760_),
    .B(_1765_),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6502_ (.A1(_1750_),
    .A2(_1757_),
    .Z(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6503_ (.A1(_1749_),
    .A2(_1758_),
    .B(_1767_),
    .ZN(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6504_ (.I(_0342_),
    .Z(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6505_ (.A1(_1769_),
    .A2(_0647_),
    .ZN(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6506_ (.A1(_1728_),
    .A2(_1770_),
    .Z(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6507_ (.I(_1771_),
    .ZN(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6508_ (.A1(_0438_),
    .A2(_1006_),
    .B1(_1023_),
    .B2(_4353_),
    .ZN(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6509_ (.A1(_1772_),
    .A2(_1773_),
    .ZN(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6510_ (.A1(_1735_),
    .A2(_1756_),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6511_ (.A1(_1735_),
    .A2(_1756_),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6512_ (.A1(_1751_),
    .A2(_1775_),
    .B(_1776_),
    .ZN(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6513_ (.A1(_0715_),
    .A2(_0961_),
    .ZN(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6514_ (.A1(\as2650.r0[2] ),
    .A2(_1015_),
    .ZN(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6515_ (.I(_1014_),
    .Z(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6516_ (.A1(_0342_),
    .A2(_1717_),
    .B1(_1780_),
    .B2(\as2650.r0[0] ),
    .ZN(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6517_ (.A1(_1718_),
    .A2(_1779_),
    .B1(_1781_),
    .B2(_1754_),
    .ZN(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6518_ (.A1(_0544_),
    .A2(_0981_),
    .ZN(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6519_ (.A1(\as2650.r0[1] ),
    .A2(_1015_),
    .ZN(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6520_ (.A1(_0442_),
    .A2(_1752_),
    .ZN(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6521_ (.A1(_1783_),
    .A2(_1784_),
    .A3(_1785_),
    .ZN(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6522_ (.A1(_1782_),
    .A2(_1786_),
    .ZN(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6523_ (.A1(_1778_),
    .A2(_1787_),
    .Z(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6524_ (.A1(_1777_),
    .A2(_1788_),
    .ZN(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6525_ (.A1(_1774_),
    .A2(_1789_),
    .ZN(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6526_ (.A1(_1766_),
    .A2(_1768_),
    .A3(_1790_),
    .Z(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6527_ (.I(_1791_),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6528_ (.A1(\as2650.r123_2[1][5] ),
    .A2(_1726_),
    .B1(_1792_),
    .B2(_1723_),
    .ZN(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6529_ (.A1(_1312_),
    .A2(_1697_),
    .ZN(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6530_ (.A1(_1793_),
    .A2(_1794_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6531_ (.A1(_1777_),
    .A2(_1788_),
    .ZN(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6532_ (.A1(_1772_),
    .A2(_1773_),
    .A3(_1789_),
    .B(_1795_),
    .ZN(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6533_ (.A1(_0519_),
    .A2(_1005_),
    .B1(_0649_),
    .B2(_0329_),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6534_ (.A1(_0443_),
    .A2(_0648_),
    .ZN(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6535_ (.A1(_1749_),
    .A2(_1798_),
    .ZN(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6536_ (.A1(_1797_),
    .A2(_1799_),
    .ZN(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6537_ (.A1(_1782_),
    .A2(_1786_),
    .ZN(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6538_ (.A1(_1778_),
    .A2(_1787_),
    .B(_1801_),
    .ZN(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6539_ (.A1(_0743_),
    .A2(_1038_),
    .Z(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6540_ (.A1(_0744_),
    .A2(_0960_),
    .B1(_1038_),
    .B2(_4316_),
    .ZN(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6541_ (.A1(_1700_),
    .A2(_1803_),
    .B(_1804_),
    .ZN(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6542_ (.A1(\as2650.r0[3] ),
    .A2(_1014_),
    .ZN(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6543_ (.A1(_0442_),
    .A2(_1717_),
    .B1(_1780_),
    .B2(\as2650.r0[1] ),
    .ZN(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6544_ (.A1(_1737_),
    .A2(_1806_),
    .B1(_1807_),
    .B2(_1783_),
    .ZN(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6545_ (.A1(\as2650.r0[5] ),
    .A2(_0980_),
    .ZN(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6546_ (.A1(_0544_),
    .A2(_1752_),
    .ZN(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6547_ (.A1(_1779_),
    .A2(_1809_),
    .A3(_1810_),
    .ZN(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6548_ (.A1(_1808_),
    .A2(_1811_),
    .Z(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6549_ (.A1(_1805_),
    .A2(_1812_),
    .Z(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6550_ (.A1(_1802_),
    .A2(_1813_),
    .Z(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6551_ (.A1(_1800_),
    .A2(_1814_),
    .Z(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6552_ (.A1(_1796_),
    .A2(_1815_),
    .ZN(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6553_ (.A1(_1771_),
    .A2(_1816_),
    .Z(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6554_ (.A1(_1768_),
    .A2(_1790_),
    .ZN(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6555_ (.A1(_1768_),
    .A2(_1790_),
    .ZN(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6556_ (.A1(_1766_),
    .A2(_1818_),
    .B(_1819_),
    .ZN(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6557_ (.A1(_1817_),
    .A2(_1820_),
    .ZN(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6558_ (.I(_1821_),
    .ZN(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6559_ (.A1(\as2650.r123_2[1][6] ),
    .A2(_1726_),
    .B1(_1822_),
    .B2(_1723_),
    .ZN(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6560_ (.A1(_1331_),
    .A2(_1696_),
    .B(_1823_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6561_ (.A1(_1817_),
    .A2(_1820_),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6562_ (.A1(_1796_),
    .A2(_1815_),
    .ZN(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6563_ (.A1(_1771_),
    .A2(_1816_),
    .B(_1825_),
    .ZN(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6564_ (.A1(_1802_),
    .A2(_1813_),
    .B1(_1814_),
    .B2(_1800_),
    .ZN(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6565_ (.A1(_1701_),
    .A2(_1803_),
    .ZN(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6566_ (.A1(_1770_),
    .A2(_1828_),
    .Z(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6567_ (.A1(_0611_),
    .A2(_1005_),
    .ZN(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6568_ (.A1(_1829_),
    .A2(_1830_),
    .Z(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6569_ (.A1(_1808_),
    .A2(_1811_),
    .B1(_1812_),
    .B2(_1805_),
    .ZN(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6570_ (.A1(_1734_),
    .A2(_1037_),
    .ZN(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6571_ (.A1(\as2650.r0[7] ),
    .A2(_0959_),
    .ZN(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6572_ (.I0(\as2650.r123[0][7] ),
    .I1(\as2650.r123_2[0][7] ),
    .S(_4108_),
    .Z(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6573_ (.A1(\as2650.r0[0] ),
    .A2(_1835_),
    .ZN(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6574_ (.A1(_1834_),
    .A2(_1836_),
    .ZN(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6575_ (.A1(_1833_),
    .A2(_1837_),
    .Z(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6576_ (.A1(\as2650.r0[4] ),
    .A2(_1014_),
    .ZN(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6577_ (.A1(_0544_),
    .A2(_1752_),
    .B1(_1780_),
    .B2(\as2650.r0[2] ),
    .ZN(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6578_ (.A1(_1753_),
    .A2(_1839_),
    .B1(_1840_),
    .B2(_1809_),
    .ZN(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6579_ (.A1(\as2650.r0[6] ),
    .A2(_0980_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6580_ (.A1(_0650_),
    .A2(_0994_),
    .ZN(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6581_ (.A1(_1806_),
    .A2(_1842_),
    .A3(_1843_),
    .ZN(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6582_ (.A1(_1841_),
    .A2(_1844_),
    .Z(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6583_ (.A1(_1838_),
    .A2(_1845_),
    .ZN(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6584_ (.A1(_1832_),
    .A2(_1846_),
    .ZN(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6585_ (.A1(_1831_),
    .A2(_1847_),
    .Z(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6586_ (.A1(_1827_),
    .A2(_1848_),
    .ZN(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6587_ (.A1(_1799_),
    .A2(_1849_),
    .Z(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6588_ (.A1(_1824_),
    .A2(_1826_),
    .A3(_1850_),
    .Z(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6589_ (.I(_1851_),
    .ZN(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6590_ (.A1(\as2650.r123_2[1][7] ),
    .A2(_1726_),
    .B1(_1852_),
    .B2(_1702_),
    .ZN(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6591_ (.A1(_1346_),
    .A2(_1696_),
    .B(_1853_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6592_ (.I(_4495_),
    .Z(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6593_ (.A1(_1046_),
    .A2(_1854_),
    .A3(_1051_),
    .ZN(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6594_ (.I(_1855_),
    .Z(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6595_ (.I(_1855_),
    .Z(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6596_ (.A1(\as2650.stack[5][0] ),
    .A2(_1857_),
    .ZN(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6597_ (.A1(_1062_),
    .A2(_1856_),
    .B(_1858_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6598_ (.A1(\as2650.stack[5][1] ),
    .A2(_1857_),
    .ZN(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6599_ (.A1(_1071_),
    .A2(_1856_),
    .B(_1859_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6600_ (.A1(\as2650.stack[5][2] ),
    .A2(_1857_),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6601_ (.A1(_1079_),
    .A2(_1856_),
    .B(_1860_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6602_ (.A1(\as2650.stack[5][3] ),
    .A2(_1857_),
    .ZN(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6603_ (.A1(_1087_),
    .A2(_1856_),
    .B(_1861_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6604_ (.I(_1855_),
    .Z(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6605_ (.I(_1855_),
    .Z(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6606_ (.A1(\as2650.stack[5][4] ),
    .A2(_1863_),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6607_ (.A1(_1093_),
    .A2(_1862_),
    .B(_1864_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6608_ (.A1(\as2650.stack[5][5] ),
    .A2(_1863_),
    .ZN(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6609_ (.A1(_1100_),
    .A2(_1862_),
    .B(_1865_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6610_ (.A1(\as2650.stack[5][6] ),
    .A2(_1863_),
    .ZN(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6611_ (.A1(_1108_),
    .A2(_1862_),
    .B(_1866_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6612_ (.A1(\as2650.stack[5][7] ),
    .A2(_1863_),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6613_ (.A1(_1115_),
    .A2(_1862_),
    .B(_1867_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6614_ (.A1(_1140_),
    .A2(_1117_),
    .ZN(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6615_ (.I(_1868_),
    .Z(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6616_ (.I(_1869_),
    .Z(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6617_ (.I(_1869_),
    .Z(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6618_ (.A1(\as2650.stack[0][8] ),
    .A2(_1871_),
    .ZN(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6619_ (.A1(_0977_),
    .A2(_1870_),
    .B(_1872_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6620_ (.I(_1868_),
    .Z(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6621_ (.A1(\as2650.stack[0][9] ),
    .A2(_1873_),
    .ZN(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6622_ (.A1(_0990_),
    .A2(_1870_),
    .B(_1874_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6623_ (.A1(\as2650.stack[0][10] ),
    .A2(_1873_),
    .ZN(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6624_ (.A1(_1001_),
    .A2(_1870_),
    .B(_1875_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6625_ (.A1(\as2650.stack[0][11] ),
    .A2(_1873_),
    .ZN(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6626_ (.A1(_1012_),
    .A2(_1870_),
    .B(_1876_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6627_ (.A1(\as2650.stack[0][12] ),
    .A2(_1873_),
    .ZN(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6628_ (.A1(_1021_),
    .A2(_1871_),
    .B(_1877_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6629_ (.A1(\as2650.stack[0][13] ),
    .A2(_1869_),
    .ZN(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6630_ (.A1(_1028_),
    .A2(_1871_),
    .B(_1878_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6631_ (.A1(\as2650.stack[0][14] ),
    .A2(_1869_),
    .ZN(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6632_ (.A1(_1043_),
    .A2(_1871_),
    .B(_1879_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6633_ (.I(\as2650.r123[3][0] ),
    .Z(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6634_ (.I(_1880_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6635_ (.I(\as2650.r123[3][1] ),
    .Z(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6636_ (.I(_1881_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6637_ (.I(\as2650.r123[3][2] ),
    .Z(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6638_ (.I(_1882_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6639_ (.I(\as2650.r123[3][3] ),
    .Z(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6640_ (.I(_1883_),
    .Z(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6641_ (.I(\as2650.r123[3][4] ),
    .Z(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6642_ (.I(_1884_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6643_ (.I(\as2650.r123[3][5] ),
    .Z(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6644_ (.I(_1885_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6645_ (.I(\as2650.r123[3][6] ),
    .Z(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6646_ (.I(_1886_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6647_ (.I(\as2650.r123[3][7] ),
    .Z(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6648_ (.I(_1887_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6649_ (.I(_1061_),
    .Z(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6650_ (.I(_0917_),
    .Z(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6651_ (.A1(_1889_),
    .A2(_1047_),
    .A3(_1051_),
    .ZN(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6652_ (.I(_1890_),
    .Z(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6653_ (.I(_1890_),
    .Z(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6654_ (.A1(\as2650.stack[3][0] ),
    .A2(_1892_),
    .ZN(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6655_ (.A1(_1888_),
    .A2(_1891_),
    .B(_1893_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6656_ (.I(_1070_),
    .Z(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6657_ (.A1(\as2650.stack[3][1] ),
    .A2(_1892_),
    .ZN(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6658_ (.A1(_1894_),
    .A2(_1891_),
    .B(_1895_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6659_ (.I(_1078_),
    .Z(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6660_ (.A1(\as2650.stack[3][2] ),
    .A2(_1892_),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6661_ (.A1(_1896_),
    .A2(_1891_),
    .B(_1897_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6662_ (.I(_1086_),
    .Z(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6663_ (.A1(\as2650.stack[3][3] ),
    .A2(_1892_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6664_ (.A1(_1898_),
    .A2(_1891_),
    .B(_1899_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6665_ (.I(_1092_),
    .Z(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6666_ (.I(_1890_),
    .Z(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6667_ (.I(_1890_),
    .Z(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6668_ (.A1(\as2650.stack[3][4] ),
    .A2(_1902_),
    .ZN(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6669_ (.A1(_1900_),
    .A2(_1901_),
    .B(_1903_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6670_ (.I(_1099_),
    .Z(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6671_ (.A1(\as2650.stack[3][5] ),
    .A2(_1902_),
    .ZN(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6672_ (.A1(_1904_),
    .A2(_1901_),
    .B(_1905_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6673_ (.I(_1107_),
    .Z(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6674_ (.A1(\as2650.stack[3][6] ),
    .A2(_1902_),
    .ZN(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6675_ (.A1(_1906_),
    .A2(_1901_),
    .B(_1907_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6676_ (.I(_1114_),
    .Z(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6677_ (.A1(\as2650.stack[3][7] ),
    .A2(_1902_),
    .ZN(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6678_ (.A1(_1908_),
    .A2(_1901_),
    .B(_1909_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6679_ (.A1(_1367_),
    .A2(_1177_),
    .ZN(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6680_ (.I(_1910_),
    .Z(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6681_ (.A1(_1693_),
    .A2(_1694_),
    .A3(_1910_),
    .ZN(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6682_ (.I(_1912_),
    .Z(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6683_ (.A1(_1217_),
    .A2(_1911_),
    .B1(_1913_),
    .B2(\as2650.r123_2[2][0] ),
    .ZN(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6684_ (.I(_1702_),
    .Z(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6685_ (.A1(_1826_),
    .A2(_1850_),
    .ZN(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6686_ (.A1(_1826_),
    .A2(_1850_),
    .ZN(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6687_ (.A1(_1824_),
    .A2(_1916_),
    .B(_1917_),
    .ZN(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6688_ (.I(_1827_),
    .ZN(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6689_ (.A1(_1919_),
    .A2(_1848_),
    .ZN(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6690_ (.A1(_1799_),
    .A2(_1849_),
    .ZN(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6691_ (.A1(_1920_),
    .A2(_1921_),
    .ZN(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6692_ (.A1(_0612_),
    .A2(_1006_),
    .A3(_1829_),
    .ZN(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6693_ (.A1(_1770_),
    .A2(_1828_),
    .B(_1923_),
    .ZN(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6694_ (.A1(_1832_),
    .A2(_1846_),
    .Z(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6695_ (.A1(_1831_),
    .A2(_1847_),
    .B(_1925_),
    .ZN(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6696_ (.A1(_4358_),
    .A2(_1835_),
    .Z(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6697_ (.A1(_1833_),
    .A2(_1837_),
    .ZN(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6698_ (.A1(_1700_),
    .A2(_1927_),
    .B(_1928_),
    .ZN(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6699_ (.A1(_1798_),
    .A2(_1929_),
    .Z(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6700_ (.A1(_0716_),
    .A2(_1004_),
    .ZN(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6701_ (.A1(_1930_),
    .A2(_1931_),
    .ZN(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6702_ (.A1(_1841_),
    .A2(_1844_),
    .ZN(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6703_ (.A1(_1838_),
    .A2(_1845_),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6704_ (.A1(_1933_),
    .A2(_1934_),
    .ZN(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6705_ (.A1(_1734_),
    .A2(_1835_),
    .ZN(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6706_ (.A1(_1769_),
    .A2(_1038_),
    .ZN(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6707_ (.A1(_1936_),
    .A2(_1937_),
    .Z(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6708_ (.A1(_0650_),
    .A2(_1780_),
    .ZN(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6709_ (.A1(_1806_),
    .A2(_1843_),
    .Z(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6710_ (.A1(_1785_),
    .A2(_1939_),
    .B1(_1940_),
    .B2(_1842_),
    .ZN(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6711_ (.A1(_0743_),
    .A2(_0993_),
    .ZN(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6712_ (.A1(_1839_),
    .A2(_1942_),
    .ZN(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6713_ (.A1(\as2650.r0[7] ),
    .A2(_0981_),
    .ZN(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6714_ (.A1(_1943_),
    .A2(_1944_),
    .Z(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6715_ (.A1(_1941_),
    .A2(_1945_),
    .Z(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6716_ (.A1(_1938_),
    .A2(_1946_),
    .Z(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6717_ (.A1(_1935_),
    .A2(_1947_),
    .Z(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6718_ (.A1(_1932_),
    .A2(_1948_),
    .Z(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6719_ (.A1(_1926_),
    .A2(_1949_),
    .Z(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6720_ (.A1(_1924_),
    .A2(_1950_),
    .Z(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6721_ (.A1(_1922_),
    .A2(_1951_),
    .Z(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6722_ (.A1(_1918_),
    .A2(_1952_),
    .Z(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6723_ (.A1(_1915_),
    .A2(_1953_),
    .ZN(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6724_ (.A1(_1914_),
    .A2(_1954_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6725_ (.A1(_1247_),
    .A2(_1911_),
    .B1(_1913_),
    .B2(\as2650.r123_2[2][1] ),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6726_ (.A1(_1922_),
    .A2(_1951_),
    .Z(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6727_ (.A1(_1918_),
    .A2(_1952_),
    .B(_1956_),
    .ZN(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6728_ (.A1(_1926_),
    .A2(_1949_),
    .Z(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6729_ (.A1(_1924_),
    .A2(_1950_),
    .B(_1958_),
    .ZN(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6730_ (.A1(_0782_),
    .A2(_1007_),
    .A3(_1930_),
    .ZN(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6731_ (.A1(_1798_),
    .A2(_1929_),
    .B(_1960_),
    .ZN(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6732_ (.A1(_1935_),
    .A2(_1947_),
    .ZN(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6733_ (.A1(_1932_),
    .A2(_1948_),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6734_ (.A1(_1962_),
    .A2(_1963_),
    .ZN(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6735_ (.A1(_1936_),
    .A2(_1937_),
    .ZN(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6736_ (.A1(_0611_),
    .A2(_0648_),
    .ZN(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6737_ (.A1(_0744_),
    .A2(_1004_),
    .ZN(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6738_ (.A1(_1965_),
    .A2(_1966_),
    .A3(_1967_),
    .Z(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6739_ (.A1(_1941_),
    .A2(_1945_),
    .ZN(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6740_ (.A1(_1938_),
    .A2(_1946_),
    .ZN(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6741_ (.A1(_1969_),
    .A2(_1970_),
    .ZN(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6742_ (.A1(_4358_),
    .A2(_0995_),
    .ZN(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6743_ (.A1(\as2650.r0[7] ),
    .A2(_1015_),
    .ZN(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6744_ (.A1(_1843_),
    .A2(_1973_),
    .ZN(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6745_ (.A1(_1939_),
    .A2(_1972_),
    .B(_1974_),
    .ZN(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6746_ (.A1(_0743_),
    .A2(_1016_),
    .ZN(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6747_ (.A1(_1810_),
    .A2(_1976_),
    .B1(_1943_),
    .B2(_1944_),
    .ZN(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6748_ (.A1(_1975_),
    .A2(_1977_),
    .Z(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6749_ (.I(_1835_),
    .Z(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6750_ (.A1(_1769_),
    .A2(_1979_),
    .B1(_1039_),
    .B2(_0444_),
    .ZN(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6751_ (.A1(_0443_),
    .A2(_1769_),
    .A3(_1979_),
    .A4(_1039_),
    .Z(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6752_ (.A1(_1980_),
    .A2(_1981_),
    .ZN(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6753_ (.A1(_1978_),
    .A2(_1982_),
    .Z(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6754_ (.A1(_1971_),
    .A2(_1983_),
    .Z(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6755_ (.A1(_1968_),
    .A2(_1984_),
    .Z(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6756_ (.A1(_1964_),
    .A2(_1985_),
    .Z(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6757_ (.A1(_1961_),
    .A2(_1986_),
    .ZN(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6758_ (.A1(_1959_),
    .A2(_1987_),
    .ZN(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6759_ (.A1(_1957_),
    .A2(_1988_),
    .Z(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6760_ (.A1(_1915_),
    .A2(_1989_),
    .ZN(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6761_ (.A1(_1955_),
    .A2(_1990_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6762_ (.A1(_1265_),
    .A2(_1911_),
    .B1(_1913_),
    .B2(\as2650.r123_2[2][2] ),
    .ZN(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6763_ (.A1(_1959_),
    .A2(_1987_),
    .Z(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6764_ (.A1(_1957_),
    .A2(_1988_),
    .B(_1992_),
    .ZN(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6765_ (.A1(_1964_),
    .A2(_1985_),
    .Z(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6766_ (.A1(_1961_),
    .A2(_1986_),
    .B(_1994_),
    .ZN(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6767_ (.A1(_0612_),
    .A2(_1023_),
    .B(_1965_),
    .ZN(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6768_ (.A1(_0644_),
    .A2(_1024_),
    .A3(_1965_),
    .ZN(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6769_ (.A1(_1996_),
    .A2(_1967_),
    .B(_1997_),
    .ZN(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6770_ (.A1(_1971_),
    .A2(_1983_),
    .ZN(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6771_ (.A1(_1968_),
    .A2(_1984_),
    .ZN(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6772_ (.A1(_1999_),
    .A2(_2000_),
    .ZN(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6773_ (.A1(_1975_),
    .A2(_1977_),
    .ZN(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6774_ (.A1(_1978_),
    .A2(_1982_),
    .ZN(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6775_ (.A1(_2002_),
    .A2(_2003_),
    .ZN(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6776_ (.I0(_1976_),
    .I1(_0744_),
    .S(_1974_),
    .Z(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6777_ (.A1(_0443_),
    .A2(_1979_),
    .ZN(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6778_ (.A1(_0545_),
    .A2(_1039_),
    .ZN(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6779_ (.A1(_2006_),
    .A2(_2007_),
    .ZN(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6780_ (.A1(_2006_),
    .A2(_2007_),
    .Z(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6781_ (.A1(_2008_),
    .A2(_2009_),
    .ZN(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6782_ (.A1(_2005_),
    .A2(_2010_),
    .ZN(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6783_ (.A1(_2004_),
    .A2(_2011_),
    .Z(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6784_ (.A1(_0715_),
    .A2(_0648_),
    .ZN(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6785_ (.A1(_1981_),
    .A2(_2013_),
    .ZN(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6786_ (.A1(_4359_),
    .A2(_1006_),
    .ZN(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6787_ (.A1(_2014_),
    .A2(_2015_),
    .Z(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6788_ (.A1(_2012_),
    .A2(_2016_),
    .Z(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6789_ (.A1(_2001_),
    .A2(_2017_),
    .Z(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6790_ (.A1(_1998_),
    .A2(_2018_),
    .ZN(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6791_ (.A1(_1995_),
    .A2(_2019_),
    .Z(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6792_ (.A1(_1993_),
    .A2(_2020_),
    .Z(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6793_ (.A1(_1915_),
    .A2(_2021_),
    .ZN(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6794_ (.A1(_1991_),
    .A2(_2022_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6795_ (.A1(_1283_),
    .A2(_1911_),
    .B1(_1913_),
    .B2(\as2650.r123_2[2][3] ),
    .ZN(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6796_ (.A1(_1995_),
    .A2(_2019_),
    .ZN(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6797_ (.A1(_1993_),
    .A2(_2020_),
    .B(_2024_),
    .ZN(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6798_ (.A1(_2001_),
    .A2(_2017_),
    .ZN(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6799_ (.A1(_1998_),
    .A2(_2018_),
    .ZN(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6800_ (.A1(_0782_),
    .A2(_1024_),
    .A3(_1981_),
    .ZN(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6801_ (.A1(_0859_),
    .A2(_1007_),
    .A3(_2014_),
    .ZN(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6802_ (.A1(_2028_),
    .A2(_2029_),
    .ZN(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6803_ (.I(_2011_),
    .ZN(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6804_ (.A1(_2004_),
    .A2(_2031_),
    .ZN(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6805_ (.A1(_2012_),
    .A2(_2016_),
    .B(_2032_),
    .ZN(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6806_ (.A1(_0745_),
    .A2(_1023_),
    .ZN(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6807_ (.A1(_2009_),
    .A2(_2034_),
    .ZN(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6808_ (.I(_1979_),
    .Z(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6809_ (.A1(_0611_),
    .A2(_2036_),
    .ZN(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6810_ (.A1(_0715_),
    .A2(_1040_),
    .ZN(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6811_ (.A1(_1973_),
    .A2(_2037_),
    .A3(_2038_),
    .ZN(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6812_ (.A1(_0793_),
    .A2(_1843_),
    .A3(_1973_),
    .B1(_2005_),
    .B2(_2010_),
    .ZN(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6813_ (.A1(_2039_),
    .A2(_2040_),
    .Z(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6814_ (.I(_2041_),
    .ZN(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6815_ (.A1(_2035_),
    .A2(_2042_),
    .Z(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6816_ (.A1(_2033_),
    .A2(_2043_),
    .ZN(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6817_ (.A1(_2030_),
    .A2(_2044_),
    .Z(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6818_ (.A1(_2026_),
    .A2(_2027_),
    .A3(_2045_),
    .Z(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6819_ (.A1(_2026_),
    .A2(_2027_),
    .B(_2045_),
    .ZN(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6820_ (.A1(_2046_),
    .A2(_2047_),
    .ZN(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6821_ (.A1(_2025_),
    .A2(_2048_),
    .ZN(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6822_ (.A1(_1915_),
    .A2(_2049_),
    .ZN(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6823_ (.A1(_2023_),
    .A2(_2050_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6824_ (.A1(_2028_),
    .A2(_2029_),
    .B(_2044_),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6825_ (.A1(_2033_),
    .A2(_2043_),
    .B(_2051_),
    .ZN(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6826_ (.A1(_2009_),
    .A2(_2034_),
    .ZN(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6827_ (.A1(_2039_),
    .A2(_2040_),
    .ZN(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6828_ (.A1(_2035_),
    .A2(_2042_),
    .B(_2054_),
    .ZN(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6829_ (.A1(_2037_),
    .A2(_2038_),
    .ZN(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6830_ (.A1(_4358_),
    .A2(_0649_),
    .Z(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6831_ (.A1(_2056_),
    .A2(_2057_),
    .ZN(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6832_ (.A1(_2037_),
    .A2(_2038_),
    .Z(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6833_ (.A1(_1973_),
    .A2(_2056_),
    .A3(_2059_),
    .ZN(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6834_ (.I(_1803_),
    .Z(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6835_ (.A1(_0716_),
    .A2(_2036_),
    .ZN(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6836_ (.A1(_2061_),
    .A2(_2062_),
    .ZN(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6837_ (.A1(_2060_),
    .A2(_2063_),
    .ZN(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6838_ (.A1(_2058_),
    .A2(_2064_),
    .Z(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6839_ (.A1(_2055_),
    .A2(_2065_),
    .Z(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6840_ (.A1(_2053_),
    .A2(_2066_),
    .ZN(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6841_ (.A1(_2052_),
    .A2(_2067_),
    .ZN(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6842_ (.A1(_1993_),
    .A2(_2020_),
    .B(_2047_),
    .C(_2024_),
    .ZN(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6843_ (.A1(_2046_),
    .A2(_2069_),
    .ZN(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6844_ (.A1(_2068_),
    .A2(_2070_),
    .Z(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6845_ (.I(_1910_),
    .Z(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6846_ (.I(_1912_),
    .Z(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6847_ (.A1(_1297_),
    .A2(_2072_),
    .B1(_2073_),
    .B2(\as2650.r123_2[2][4] ),
    .ZN(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6848_ (.A1(_1298_),
    .A2(_2071_),
    .B(_2074_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6849_ (.A1(_1312_),
    .A2(_2072_),
    .B1(_2073_),
    .B2(\as2650.r123_2[2][5] ),
    .ZN(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6850_ (.A1(_2055_),
    .A2(_2065_),
    .ZN(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6851_ (.A1(_2053_),
    .A2(_2066_),
    .ZN(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6852_ (.A1(_2076_),
    .A2(_2077_),
    .ZN(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6853_ (.I(_2078_),
    .ZN(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6854_ (.A1(_2060_),
    .A2(_2063_),
    .ZN(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6855_ (.A1(_2058_),
    .A2(_2064_),
    .B(_2080_),
    .ZN(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6856_ (.I(_2036_),
    .Z(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6857_ (.A1(_0822_),
    .A2(_2082_),
    .B1(_1040_),
    .B2(_0859_),
    .ZN(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6858_ (.A1(_0859_),
    .A2(_2036_),
    .A3(_2061_),
    .Z(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6859_ (.A1(_2083_),
    .A2(_2084_),
    .ZN(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6860_ (.A1(_0782_),
    .A2(_2082_),
    .A3(_2061_),
    .ZN(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6861_ (.I0(_0860_),
    .I1(_2085_),
    .S(_2086_),
    .Z(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6862_ (.A1(_2056_),
    .A2(_2057_),
    .B1(_2081_),
    .B2(_2087_),
    .ZN(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6863_ (.A1(_2081_),
    .A2(_2087_),
    .B(_2088_),
    .ZN(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6864_ (.A1(_2046_),
    .A2(_2068_),
    .A3(_2069_),
    .B1(_2052_),
    .B2(_2067_),
    .ZN(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6865_ (.A1(_2079_),
    .A2(_2089_),
    .A3(_2090_),
    .Z(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6866_ (.A1(_1703_),
    .A2(_2091_),
    .ZN(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6867_ (.A1(_2075_),
    .A2(_2092_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6868_ (.A1(_1332_),
    .A2(_2072_),
    .B1(_2073_),
    .B2(\as2650.r123_2[2][6] ),
    .ZN(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6869_ (.A1(_2079_),
    .A2(_2089_),
    .ZN(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6870_ (.A1(_2079_),
    .A2(_2089_),
    .ZN(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6871_ (.A1(_2094_),
    .A2(_2090_),
    .B(_2095_),
    .ZN(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6872_ (.A1(_0909_),
    .A2(_2082_),
    .ZN(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _6873_ (.A1(_2061_),
    .A2(_2097_),
    .B1(_2086_),
    .B2(_0909_),
    .ZN(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6874_ (.A1(_2088_),
    .A2(_2098_),
    .Z(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6875_ (.A1(_2096_),
    .A2(_2099_),
    .Z(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6876_ (.A1(_1703_),
    .A2(_2100_),
    .ZN(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6877_ (.A1(_2093_),
    .A2(_2101_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6878_ (.I(_2072_),
    .ZN(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6879_ (.I(_2088_),
    .ZN(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6880_ (.A1(_2096_),
    .A2(_2099_),
    .ZN(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6881_ (.A1(_2103_),
    .A2(_2098_),
    .B(_2104_),
    .C(_2084_),
    .ZN(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6882_ (.A1(\as2650.r123_2[2][7] ),
    .A2(_2073_),
    .ZN(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6883_ (.A1(_1346_),
    .A2(_2102_),
    .B1(_2105_),
    .B2(_1298_),
    .C(_2106_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6884_ (.A1(_1045_),
    .A2(_1854_),
    .A3(_1118_),
    .ZN(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6885_ (.I(_2107_),
    .Z(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6886_ (.I(_2107_),
    .Z(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6887_ (.A1(\as2650.stack[4][0] ),
    .A2(_2109_),
    .ZN(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6888_ (.A1(_1888_),
    .A2(_2108_),
    .B(_2110_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6889_ (.A1(\as2650.stack[4][1] ),
    .A2(_2109_),
    .ZN(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6890_ (.A1(_1894_),
    .A2(_2108_),
    .B(_2111_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6891_ (.A1(\as2650.stack[4][2] ),
    .A2(_2109_),
    .ZN(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6892_ (.A1(_1896_),
    .A2(_2108_),
    .B(_2112_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6893_ (.A1(\as2650.stack[4][3] ),
    .A2(_2109_),
    .ZN(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6894_ (.A1(_1898_),
    .A2(_2108_),
    .B(_2113_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6895_ (.I(_2107_),
    .Z(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6896_ (.I(_2107_),
    .Z(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6897_ (.A1(\as2650.stack[4][4] ),
    .A2(_2115_),
    .ZN(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6898_ (.A1(_1900_),
    .A2(_2114_),
    .B(_2116_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6899_ (.A1(\as2650.stack[4][5] ),
    .A2(_2115_),
    .ZN(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6900_ (.A1(_1904_),
    .A2(_2114_),
    .B(_2117_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6901_ (.A1(\as2650.stack[4][6] ),
    .A2(_2115_),
    .ZN(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6902_ (.A1(_1906_),
    .A2(_2114_),
    .B(_2118_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6903_ (.A1(\as2650.stack[4][7] ),
    .A2(_2115_),
    .ZN(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6904_ (.A1(_1908_),
    .A2(_2114_),
    .B(_2119_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6905_ (.I(_1203_),
    .Z(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6906_ (.I(_4235_),
    .Z(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6907_ (.I(\as2650.cycle[6] ),
    .Z(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6908_ (.I(_4239_),
    .Z(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6909_ (.A1(_2122_),
    .A2(_2123_),
    .A3(_4252_),
    .ZN(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6910_ (.A1(_2121_),
    .A2(_2124_),
    .ZN(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6911_ (.A1(_4425_),
    .A2(_2125_),
    .ZN(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6912_ (.I(_2126_),
    .Z(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6913_ (.A1(_4190_),
    .A2(_0949_),
    .ZN(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6914_ (.A1(_0405_),
    .A2(_2128_),
    .ZN(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6915_ (.A1(_2129_),
    .A2(_4195_),
    .ZN(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6916_ (.A1(_2121_),
    .A2(_2123_),
    .A3(_1460_),
    .ZN(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6917_ (.A1(_0928_),
    .A2(_2130_),
    .A3(_2131_),
    .Z(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6918_ (.A1(_1486_),
    .A2(_2127_),
    .A3(_2132_),
    .ZN(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6919_ (.I(_4425_),
    .Z(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6920_ (.I(_2134_),
    .Z(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6921_ (.I(_4195_),
    .Z(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6922_ (.A1(_1682_),
    .A2(_2136_),
    .ZN(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6923_ (.A1(_0970_),
    .A2(_2137_),
    .B(_1660_),
    .ZN(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _6924_ (.A1(_1512_),
    .A2(_1394_),
    .A3(_2135_),
    .B1(_1675_),
    .B2(_2138_),
    .ZN(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6925_ (.A1(_4210_),
    .A2(_1661_),
    .ZN(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6926_ (.I(_2140_),
    .Z(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6927_ (.I(_0928_),
    .Z(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6928_ (.A1(_1442_),
    .A2(_2142_),
    .ZN(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6929_ (.A1(_1372_),
    .A2(_2140_),
    .ZN(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6930_ (.I(_2128_),
    .Z(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6931_ (.A1(_0943_),
    .A2(_2145_),
    .ZN(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6932_ (.A1(_2141_),
    .A2(_1452_),
    .A3(_2143_),
    .B1(_2144_),
    .B2(_2146_),
    .ZN(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6933_ (.A1(_1662_),
    .A2(_1674_),
    .ZN(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6934_ (.A1(_0945_),
    .A2(_2147_),
    .A3(_2148_),
    .ZN(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6935_ (.I(_0948_),
    .Z(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6936_ (.A1(_1188_),
    .A2(_2150_),
    .B(_0950_),
    .C(_4421_),
    .ZN(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6937_ (.A1(_2121_),
    .A2(_2123_),
    .A3(_1460_),
    .ZN(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6938_ (.A1(_2122_),
    .A2(_2152_),
    .ZN(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6939_ (.A1(_1511_),
    .A2(_2142_),
    .B(_1671_),
    .ZN(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6940_ (.A1(_1476_),
    .A2(_2153_),
    .B(_2154_),
    .ZN(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6941_ (.I(_2155_),
    .ZN(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6942_ (.A1(_1664_),
    .A2(_1463_),
    .A3(_2151_),
    .A4(_2156_),
    .ZN(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _6943_ (.A1(_2133_),
    .A2(_2139_),
    .A3(_2149_),
    .A4(_2157_),
    .ZN(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6944_ (.I(_2158_),
    .Z(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6945_ (.I(\as2650.addr_buff[0] ),
    .Z(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6946_ (.I(_2160_),
    .Z(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6947_ (.I(_2161_),
    .Z(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6948_ (.I(_2158_),
    .Z(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6949_ (.A1(_2162_),
    .A2(_2163_),
    .ZN(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6950_ (.A1(_2120_),
    .A2(_2159_),
    .B(_2164_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6951_ (.I(\as2650.addr_buff[1] ),
    .Z(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6952_ (.A1(_2165_),
    .A2(_2163_),
    .ZN(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6953_ (.A1(_1236_),
    .A2(_2159_),
    .B(_2166_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6954_ (.I(_1609_),
    .Z(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6955_ (.I(\as2650.addr_buff[2] ),
    .Z(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6956_ (.I(_2168_),
    .Z(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6957_ (.A1(_2169_),
    .A2(_2163_),
    .ZN(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6958_ (.A1(_2167_),
    .A2(_2159_),
    .B(_2170_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6959_ (.I(_1556_),
    .Z(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6960_ (.I(\as2650.addr_buff[3] ),
    .Z(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6961_ (.I(_2172_),
    .Z(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6962_ (.I(_2158_),
    .Z(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6963_ (.I0(_2171_),
    .I1(_2173_),
    .S(_2174_),
    .Z(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6964_ (.I(_2175_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6965_ (.I(_0677_),
    .Z(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6966_ (.I(\as2650.addr_buff[4] ),
    .Z(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6967_ (.I0(_2176_),
    .I1(_2177_),
    .S(_2174_),
    .Z(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6968_ (.I(_2178_),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6969_ (.I(_1585_),
    .Z(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6970_ (.I(_4244_),
    .Z(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6971_ (.A1(_2180_),
    .A2(_2174_),
    .ZN(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6972_ (.A1(_2179_),
    .A2(_2159_),
    .B(_2181_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6973_ (.I(_4243_),
    .Z(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6974_ (.I0(_1689_),
    .I1(_2182_),
    .S(_2158_),
    .Z(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6975_ (.I(_2183_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6976_ (.I(_1581_),
    .Z(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6977_ (.I(_2184_),
    .Z(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6978_ (.I(_2185_),
    .Z(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6979_ (.I(_4427_),
    .Z(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6980_ (.A1(_2187_),
    .A2(_2174_),
    .ZN(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6981_ (.A1(_2186_),
    .A2(_2163_),
    .B(_2188_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6982_ (.I(net24),
    .ZN(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6983_ (.I(_1436_),
    .Z(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6984_ (.I(_1206_),
    .Z(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6985_ (.I(_1362_),
    .Z(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6986_ (.A1(_2191_),
    .A2(_2192_),
    .ZN(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6987_ (.A1(_0969_),
    .A2(_2193_),
    .ZN(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6988_ (.I(_2194_),
    .Z(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6989_ (.A1(_2190_),
    .A2(_2195_),
    .ZN(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6990_ (.I(_2130_),
    .Z(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6991_ (.I(_2197_),
    .Z(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6992_ (.I(_4114_),
    .Z(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6993_ (.A1(_0334_),
    .A2(_1381_),
    .A3(_2143_),
    .Z(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6994_ (.A1(_2199_),
    .A2(_2200_),
    .ZN(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6995_ (.I(_4200_),
    .Z(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6996_ (.A1(_1435_),
    .A2(_1466_),
    .A3(_2202_),
    .ZN(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6997_ (.A1(_2201_),
    .A2(_2203_),
    .ZN(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6998_ (.A1(_2142_),
    .A2(_1453_),
    .B1(_2196_),
    .B2(_2198_),
    .C(_2204_),
    .ZN(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6999_ (.I(_2129_),
    .Z(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7000_ (.A1(_2206_),
    .A2(_1485_),
    .ZN(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _7001_ (.I(_2207_),
    .ZN(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7002_ (.I(_1475_),
    .Z(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7003_ (.A1(_2209_),
    .A2(_2192_),
    .ZN(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7004_ (.A1(_1324_),
    .A2(_1363_),
    .ZN(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7005_ (.A1(_1446_),
    .A2(_1675_),
    .A3(_2210_),
    .A4(_2211_),
    .ZN(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _7006_ (.A1(_4202_),
    .A2(_1463_),
    .A3(_2208_),
    .A4(_2212_),
    .ZN(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7007_ (.A1(_2205_),
    .A2(_2213_),
    .ZN(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7008_ (.I(_1513_),
    .Z(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7009_ (.I(_2136_),
    .Z(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7010_ (.I(_2216_),
    .Z(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7011_ (.A1(_4193_),
    .A2(_4250_),
    .A3(_0928_),
    .ZN(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7012_ (.A1(_2215_),
    .A2(_2217_),
    .B(_2218_),
    .C(_2214_),
    .ZN(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7013_ (.A1(_2189_),
    .A2(_2214_),
    .B(_2219_),
    .C(_1644_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7014_ (.I(_2199_),
    .Z(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7015_ (.I(_2191_),
    .Z(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7016_ (.I(_2221_),
    .Z(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7017_ (.I(_2222_),
    .Z(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7018_ (.I(_1670_),
    .Z(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7019_ (.I(_2224_),
    .Z(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7020_ (.I(_1638_),
    .Z(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7021_ (.A1(_2202_),
    .A2(_2226_),
    .ZN(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _7022_ (.A1(_2220_),
    .A2(_2223_),
    .A3(_2225_),
    .A4(_2227_),
    .ZN(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7023_ (.A1(net22),
    .A2(_2228_),
    .ZN(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7024_ (.A1(_4141_),
    .A2(_2228_),
    .B(_2229_),
    .C(_1644_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7025_ (.I(_1424_),
    .Z(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7026_ (.I(_2230_),
    .Z(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7027_ (.A1(_0404_),
    .A2(_4123_),
    .ZN(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7028_ (.I(_2232_),
    .Z(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7029_ (.A1(_1206_),
    .A2(_1389_),
    .ZN(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7030_ (.I(_2234_),
    .Z(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7031_ (.I(_2206_),
    .Z(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7032_ (.A1(_1459_),
    .A2(_2236_),
    .B(_1373_),
    .ZN(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _7033_ (.A1(_2233_),
    .A2(_2235_),
    .B1(_2237_),
    .B2(_1437_),
    .ZN(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7034_ (.I(_4410_),
    .Z(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7035_ (.A1(_2239_),
    .A2(_2225_),
    .B(_1474_),
    .ZN(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7036_ (.A1(_2209_),
    .A2(_1422_),
    .ZN(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7037_ (.I(_1461_),
    .Z(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7038_ (.A1(_1523_),
    .A2(_2242_),
    .ZN(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7039_ (.I(_2243_),
    .Z(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7040_ (.I(_2244_),
    .Z(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7041_ (.A1(_2202_),
    .A2(_2241_),
    .A3(_2245_),
    .B1(_1574_),
    .B2(_1459_),
    .ZN(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7042_ (.A1(_2240_),
    .A2(_2246_),
    .ZN(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7043_ (.A1(_1385_),
    .A2(_2238_),
    .A3(_2247_),
    .ZN(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7044_ (.A1(_2238_),
    .A2(_2247_),
    .ZN(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7045_ (.A1(net23),
    .A2(_2249_),
    .ZN(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7046_ (.A1(_2231_),
    .A2(_2248_),
    .A3(_2250_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7047_ (.A1(_4224_),
    .A2(_4169_),
    .ZN(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7048_ (.A1(_4185_),
    .A2(_1519_),
    .A3(_2224_),
    .ZN(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7049_ (.A1(_1400_),
    .A2(_4158_),
    .A3(_1353_),
    .ZN(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7050_ (.A1(_2253_),
    .A2(_1404_),
    .B(_0944_),
    .ZN(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7051_ (.A1(_2252_),
    .A2(_2254_),
    .ZN(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7052_ (.A1(_1379_),
    .A2(_1670_),
    .ZN(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7053_ (.A1(_1359_),
    .A2(_2256_),
    .ZN(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7054_ (.A1(_2251_),
    .A2(_2255_),
    .A3(_2257_),
    .ZN(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7055_ (.I(_1441_),
    .Z(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7056_ (.A1(_4251_),
    .A2(_2224_),
    .ZN(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7057_ (.A1(_4257_),
    .A2(_0334_),
    .B(_1349_),
    .ZN(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7058_ (.A1(_4222_),
    .A2(_2259_),
    .A3(_2260_),
    .A4(_2261_),
    .ZN(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7059_ (.A1(_1033_),
    .A2(_2262_),
    .ZN(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7060_ (.I(_0929_),
    .Z(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7061_ (.A1(_4126_),
    .A2(_1379_),
    .A3(_1364_),
    .ZN(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7062_ (.A1(_2232_),
    .A2(_2265_),
    .ZN(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7063_ (.A1(_1447_),
    .A2(_2218_),
    .ZN(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7064_ (.A1(_2266_),
    .A2(_2267_),
    .ZN(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7065_ (.A1(_2233_),
    .A2(_2234_),
    .ZN(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7066_ (.A1(_4227_),
    .A2(_4199_),
    .ZN(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7067_ (.A1(_2270_),
    .A2(_2233_),
    .ZN(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7068_ (.A1(_4226_),
    .A2(_4504_),
    .A3(_0655_),
    .ZN(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7069_ (.I(_2272_),
    .Z(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7070_ (.A1(_4514_),
    .A2(_2273_),
    .B(_1386_),
    .ZN(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7071_ (.A1(_1671_),
    .A2(_2269_),
    .A3(_2271_),
    .A4(_2274_),
    .ZN(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7072_ (.A1(_1476_),
    .A2(_2264_),
    .B(_2268_),
    .C(_2275_),
    .ZN(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7073_ (.A1(_2224_),
    .A2(_2149_),
    .B(_2276_),
    .ZN(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7074_ (.A1(_2258_),
    .A2(_2263_),
    .A3(_2277_),
    .ZN(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7075_ (.A1(_2126_),
    .A2(_2132_),
    .ZN(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7076_ (.A1(_1450_),
    .A2(_2242_),
    .ZN(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7077_ (.I(_1384_),
    .Z(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7078_ (.I(_0405_),
    .Z(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7079_ (.I(_4194_),
    .Z(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7080_ (.A1(_2282_),
    .A2(_2283_),
    .ZN(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7081_ (.A1(_2281_),
    .A2(_2284_),
    .B(_2132_),
    .ZN(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _7082_ (.A1(_1252_),
    .A2(_2279_),
    .A3(_2280_),
    .A4(_2285_),
    .ZN(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7083_ (.A1(_4234_),
    .A2(_1459_),
    .A3(_0939_),
    .ZN(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7084_ (.I(_4115_),
    .Z(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7085_ (.A1(_1523_),
    .A2(_1373_),
    .B(_2288_),
    .ZN(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _7086_ (.A1(_2208_),
    .A2(_2286_),
    .A3(_2287_),
    .A4(_2289_),
    .ZN(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7087_ (.A1(_2278_),
    .A2(_2290_),
    .ZN(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7088_ (.A1(_2191_),
    .A2(_0923_),
    .ZN(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7089_ (.A1(_0663_),
    .A2(_0761_),
    .Z(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7090_ (.A1(_4399_),
    .A2(_0361_),
    .A3(_0463_),
    .A4(_0560_),
    .ZN(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7091_ (.A1(_0673_),
    .A2(_2294_),
    .Z(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _7092_ (.A1(_2293_),
    .A2(_0829_),
    .A3(_0898_),
    .A4(_2295_),
    .Z(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7093_ (.A1(_4512_),
    .A2(_1356_),
    .B(_1357_),
    .ZN(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7094_ (.A1(_4183_),
    .A2(_2296_),
    .B(_2297_),
    .ZN(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7095_ (.A1(_4206_),
    .A2(_2298_),
    .ZN(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7096_ (.A1(_4133_),
    .A2(_4145_),
    .A3(_1353_),
    .ZN(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7097_ (.A1(_2259_),
    .A2(_2300_),
    .ZN(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7098_ (.A1(_4224_),
    .A2(_2301_),
    .ZN(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7099_ (.A1(_2292_),
    .A2(_2299_),
    .B(_2302_),
    .ZN(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7100_ (.A1(_2291_),
    .A2(_2303_),
    .ZN(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7101_ (.I(_2304_),
    .Z(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7102_ (.I(_2305_),
    .Z(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7103_ (.I(_2306_),
    .Z(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7104_ (.I(_2242_),
    .Z(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7105_ (.I(_2308_),
    .Z(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7106_ (.I(_1056_),
    .Z(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7107_ (.I(_2310_),
    .Z(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7108_ (.A1(_2221_),
    .A2(_1188_),
    .ZN(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7109_ (.I(_2312_),
    .Z(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7110_ (.A1(_0938_),
    .A2(_1455_),
    .ZN(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7111_ (.I(_2314_),
    .Z(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7112_ (.A1(_2313_),
    .A2(_2315_),
    .ZN(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7113_ (.I(_1572_),
    .Z(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7114_ (.A1(_2311_),
    .A2(_2316_),
    .B(_2317_),
    .ZN(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7115_ (.I(net54),
    .ZN(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7116_ (.I(_1543_),
    .Z(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7117_ (.I(_2320_),
    .Z(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7118_ (.I(_2321_),
    .Z(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7119_ (.I(_0902_),
    .Z(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7120_ (.I(_2323_),
    .Z(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7121_ (.A1(_2310_),
    .A2(_1549_),
    .Z(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7122_ (.A1(_2324_),
    .A2(_2325_),
    .ZN(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7123_ (.I(_0939_),
    .Z(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7124_ (.A1(_2137_),
    .A2(_2327_),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7125_ (.I(_2328_),
    .Z(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7126_ (.A1(_2319_),
    .A2(_2322_),
    .B(_2326_),
    .C(_2329_),
    .ZN(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7127_ (.I(_4426_),
    .ZN(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7128_ (.I(_2331_),
    .Z(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7129_ (.I(_2129_),
    .Z(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7130_ (.I(_2333_),
    .Z(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7131_ (.I(_2334_),
    .Z(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7132_ (.A1(_1549_),
    .A2(_2335_),
    .ZN(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7133_ (.I(net54),
    .Z(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7134_ (.I(_4256_),
    .Z(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7135_ (.I(_2338_),
    .Z(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7136_ (.I(_2206_),
    .Z(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7137_ (.A1(_2332_),
    .A2(_2340_),
    .ZN(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7138_ (.A1(_2337_),
    .A2(_2341_),
    .ZN(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7139_ (.A1(_2337_),
    .A2(_2339_),
    .B(_2342_),
    .ZN(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7140_ (.I(_1663_),
    .Z(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7141_ (.A1(_2216_),
    .A2(_2344_),
    .ZN(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7142_ (.I(_2345_),
    .Z(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7143_ (.A1(_2332_),
    .A2(_2336_),
    .B(_2343_),
    .C(_2346_),
    .ZN(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7144_ (.I(_2313_),
    .Z(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7145_ (.A1(_2330_),
    .A2(_2347_),
    .B(_2348_),
    .ZN(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7146_ (.I(_2131_),
    .Z(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7147_ (.I(_2350_),
    .ZN(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7148_ (.I(_2351_),
    .Z(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7149_ (.I(_2126_),
    .Z(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7150_ (.I(_2353_),
    .Z(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7151_ (.A1(_4447_),
    .A2(_4459_),
    .ZN(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7152_ (.A1(_1549_),
    .A2(_2355_),
    .Z(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7153_ (.I(_4246_),
    .Z(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7154_ (.I(_2357_),
    .Z(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7155_ (.A1(_2358_),
    .A2(_4438_),
    .ZN(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7156_ (.A1(_2120_),
    .A2(_2359_),
    .Z(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7157_ (.I(_2134_),
    .Z(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7158_ (.I(_2361_),
    .Z(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7159_ (.A1(_2354_),
    .A2(_2356_),
    .B1(_2360_),
    .B2(_2362_),
    .ZN(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7160_ (.A1(_4240_),
    .A2(_2282_),
    .ZN(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7161_ (.I(_2364_),
    .Z(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7162_ (.I(_2122_),
    .Z(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7163_ (.A1(_2366_),
    .A2(_2131_),
    .ZN(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7164_ (.I(_2367_),
    .Z(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7165_ (.A1(_2337_),
    .A2(_2365_),
    .B1(_2368_),
    .B2(_2325_),
    .ZN(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7166_ (.I(_1487_),
    .Z(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7167_ (.A1(_2352_),
    .A2(_2363_),
    .B(_2369_),
    .C(_2370_),
    .ZN(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7168_ (.A1(_2318_),
    .A2(_2349_),
    .B(_2371_),
    .ZN(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7169_ (.I(_1446_),
    .Z(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7170_ (.I(_2308_),
    .Z(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7171_ (.A1(_2373_),
    .A2(_2374_),
    .ZN(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7172_ (.A1(_2309_),
    .A2(_2372_),
    .B1(_2375_),
    .B2(_2311_),
    .ZN(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7173_ (.I(_2304_),
    .Z(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7174_ (.A1(_2337_),
    .A2(_2377_),
    .B(_1425_),
    .ZN(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7175_ (.A1(_2307_),
    .A2(_2376_),
    .B(_2378_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7176_ (.I(_2305_),
    .Z(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7177_ (.I(_1066_),
    .Z(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7178_ (.A1(_2281_),
    .A2(_2282_),
    .ZN(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7179_ (.I(_2381_),
    .Z(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7180_ (.A1(_1564_),
    .A2(_2382_),
    .ZN(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7181_ (.I(_2383_),
    .Z(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7182_ (.I(_1451_),
    .Z(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7183_ (.I(_2385_),
    .Z(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7184_ (.I(_4447_),
    .Z(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7185_ (.I(_2353_),
    .Z(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7186_ (.I(_4446_),
    .Z(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7187_ (.A1(_4386_),
    .A2(_4458_),
    .ZN(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7188_ (.A1(_0352_),
    .A2(_0320_),
    .A3(_2390_),
    .Z(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7189_ (.A1(_2389_),
    .A2(_2391_),
    .ZN(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7190_ (.A1(_1551_),
    .A2(_2387_),
    .B(_2388_),
    .C(_2392_),
    .ZN(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7191_ (.I(_4428_),
    .Z(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7192_ (.I(_2394_),
    .Z(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7193_ (.A1(_1203_),
    .A2(_4437_),
    .Z(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7194_ (.A1(_0351_),
    .A2(_0328_),
    .A3(_2396_),
    .Z(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7195_ (.A1(_2395_),
    .A2(_2397_),
    .ZN(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7196_ (.I(_2134_),
    .Z(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7197_ (.A1(_1551_),
    .A2(_2395_),
    .B(_2398_),
    .C(_2399_),
    .ZN(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7198_ (.A1(_2393_),
    .A2(_2400_),
    .B(_2352_),
    .ZN(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7199_ (.I(_2124_),
    .Z(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7200_ (.I(net29),
    .Z(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7201_ (.A1(_2403_),
    .A2(_2319_),
    .Z(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7202_ (.I(_2367_),
    .Z(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7203_ (.A1(\as2650.pc[1] ),
    .A2(net7),
    .Z(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7204_ (.A1(_1055_),
    .A2(_4386_),
    .B(_2406_),
    .ZN(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _7205_ (.A1(_2310_),
    .A2(_1550_),
    .A3(_2406_),
    .Z(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7206_ (.A1(_2405_),
    .A2(_2407_),
    .A3(_2408_),
    .ZN(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7207_ (.A1(_2402_),
    .A2(_2404_),
    .B(_2409_),
    .ZN(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7208_ (.I(_4410_),
    .Z(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7209_ (.I(_1658_),
    .Z(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7210_ (.A1(_4427_),
    .A2(_2334_),
    .ZN(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7211_ (.A1(_0408_),
    .A2(_2404_),
    .ZN(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7212_ (.A1(_2403_),
    .A2(_2341_),
    .B1(_2413_),
    .B2(_0353_),
    .C(_2414_),
    .ZN(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _7213_ (.A1(_2412_),
    .A2(_1664_),
    .A3(_2415_),
    .Z(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7214_ (.A1(_0930_),
    .A2(_4195_),
    .ZN(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7215_ (.I(_2417_),
    .Z(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7216_ (.A1(_0970_),
    .A2(_2418_),
    .ZN(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7217_ (.I(_0932_),
    .Z(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7218_ (.A1(_2420_),
    .A2(_1663_),
    .ZN(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7219_ (.A1(_1465_),
    .A2(_2421_),
    .ZN(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7220_ (.I(_2422_),
    .Z(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7221_ (.A1(_1055_),
    .A2(net6),
    .ZN(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7222_ (.A1(_2424_),
    .A2(_2406_),
    .Z(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7223_ (.I(_1620_),
    .Z(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7224_ (.A1(_2403_),
    .A2(_2426_),
    .ZN(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7225_ (.A1(_2323_),
    .A2(_2425_),
    .B(_2427_),
    .ZN(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7226_ (.A1(_2380_),
    .A2(_2419_),
    .B1(_2423_),
    .B2(_2428_),
    .C(_1676_),
    .ZN(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7227_ (.A1(_1068_),
    .A2(_2411_),
    .B1(_2416_),
    .B2(_2429_),
    .ZN(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7228_ (.A1(_2386_),
    .A2(_2401_),
    .A3(_2410_),
    .B(_2430_),
    .ZN(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7229_ (.A1(_2374_),
    .A2(_2431_),
    .ZN(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7230_ (.A1(_2380_),
    .A2(_2384_),
    .B(_2432_),
    .ZN(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7231_ (.I(_2305_),
    .Z(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7232_ (.A1(_2403_),
    .A2(_2434_),
    .ZN(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7233_ (.I(_1693_),
    .Z(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7234_ (.I(_2436_),
    .Z(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7235_ (.A1(_2379_),
    .A2(_2433_),
    .B(_2435_),
    .C(_2437_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7236_ (.I(_1380_),
    .Z(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7237_ (.I(_1487_),
    .Z(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7238_ (.I(net7),
    .Z(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7239_ (.A1(_2440_),
    .A2(_0319_),
    .ZN(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7240_ (.A1(_0350_),
    .A2(_0319_),
    .ZN(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7241_ (.A1(_2390_),
    .A2(_2441_),
    .B(_2442_),
    .ZN(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7242_ (.A1(_0455_),
    .A2(_0485_),
    .Z(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7243_ (.A1(_2443_),
    .A2(_2444_),
    .B(_4278_),
    .ZN(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7244_ (.A1(_2443_),
    .A2(_2444_),
    .B(_2445_),
    .ZN(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7245_ (.A1(_1553_),
    .A2(_2389_),
    .B(_2127_),
    .C(_2446_),
    .ZN(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7246_ (.A1(_2440_),
    .A2(_0327_),
    .ZN(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7247_ (.A1(_2440_),
    .A2(_0327_),
    .ZN(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7248_ (.A1(_2448_),
    .A2(_2396_),
    .B(_2449_),
    .ZN(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7249_ (.A1(_0454_),
    .A2(_0475_),
    .Z(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7250_ (.A1(_0456_),
    .A2(_0476_),
    .ZN(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7251_ (.A1(_2451_),
    .A2(_2452_),
    .ZN(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7252_ (.A1(_2450_),
    .A2(_2453_),
    .B(_2357_),
    .ZN(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7253_ (.A1(_2450_),
    .A2(_2453_),
    .B(_2454_),
    .ZN(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7254_ (.A1(_1552_),
    .A2(_2394_),
    .B(_2455_),
    .C(_2135_),
    .ZN(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7255_ (.A1(_2447_),
    .A2(_2456_),
    .ZN(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7256_ (.A1(_2350_),
    .A2(_2457_),
    .ZN(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7257_ (.A1(\as2650.pc[2] ),
    .A2(net8),
    .Z(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7258_ (.A1(\as2650.pc[1] ),
    .A2(_0349_),
    .ZN(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7259_ (.A1(_2460_),
    .A2(_2407_),
    .ZN(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7260_ (.A1(_2459_),
    .A2(_2461_),
    .ZN(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7261_ (.A1(_1073_),
    .A2(_2167_),
    .Z(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7262_ (.A1(_2460_),
    .A2(_2407_),
    .A3(_2463_),
    .ZN(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7263_ (.A1(_2405_),
    .A2(_2462_),
    .A3(_2464_),
    .ZN(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7264_ (.I(_2364_),
    .Z(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7265_ (.I(net30),
    .Z(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7266_ (.A1(net29),
    .A2(net54),
    .ZN(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7267_ (.A1(_2467_),
    .A2(_2468_),
    .ZN(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7268_ (.A1(_2466_),
    .A2(_2469_),
    .ZN(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7269_ (.A1(_2439_),
    .A2(_2458_),
    .A3(_2465_),
    .A4(_2470_),
    .ZN(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7270_ (.I(_2341_),
    .Z(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7271_ (.A1(_2331_),
    .A2(_0935_),
    .ZN(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7272_ (.I(_2473_),
    .Z(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7273_ (.I(_0951_),
    .Z(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7274_ (.I(_2475_),
    .Z(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7275_ (.A1(_2476_),
    .A2(_2469_),
    .ZN(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7276_ (.A1(_2167_),
    .A2(_2474_),
    .B(_2477_),
    .ZN(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7277_ (.A1(_2467_),
    .A2(_2472_),
    .B(_2346_),
    .C(_2478_),
    .ZN(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7278_ (.A1(_1066_),
    .A2(_0349_),
    .ZN(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7279_ (.A1(_2424_),
    .A2(_2480_),
    .B(_2460_),
    .ZN(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7280_ (.A1(_2463_),
    .A2(_2481_),
    .Z(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7281_ (.A1(_2467_),
    .A2(_2426_),
    .ZN(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7282_ (.A1(_2323_),
    .A2(_2482_),
    .B(_2483_),
    .ZN(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7283_ (.A1(_1075_),
    .A2(_2419_),
    .B1(_2422_),
    .B2(_2484_),
    .C(_1675_),
    .ZN(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7284_ (.A1(_1395_),
    .A2(_2479_),
    .B(_2485_),
    .ZN(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7285_ (.A1(_1076_),
    .A2(_2438_),
    .B(_2471_),
    .C(_2486_),
    .ZN(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7286_ (.A1(_2308_),
    .A2(_2487_),
    .ZN(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7287_ (.A1(_1076_),
    .A2(_2384_),
    .B(_2488_),
    .ZN(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7288_ (.A1(_2467_),
    .A2(_2434_),
    .ZN(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7289_ (.A1(_2379_),
    .A2(_2489_),
    .B(_2490_),
    .C(_2437_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7290_ (.I(\as2650.pc[3] ),
    .Z(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7291_ (.I(_2491_),
    .Z(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7292_ (.I(_2383_),
    .Z(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7293_ (.A1(net30),
    .A2(net29),
    .A3(net54),
    .ZN(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7294_ (.A1(net53),
    .A2(_2494_),
    .Z(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7295_ (.A1(_2365_),
    .A2(_2495_),
    .ZN(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _7296_ (.A1(_2121_),
    .A2(_2366_),
    .A3(_2123_),
    .A4(_1460_),
    .ZN(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7297_ (.I(_4278_),
    .Z(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7298_ (.A1(_0479_),
    .A2(_0484_),
    .B(_1609_),
    .ZN(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7299_ (.A1(_1609_),
    .A2(_0479_),
    .A3(_0484_),
    .ZN(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7300_ (.A1(_2443_),
    .A2(_2499_),
    .B(_2500_),
    .ZN(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7301_ (.A1(_0556_),
    .A2(_1271_),
    .A3(_2501_),
    .Z(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7302_ (.A1(_1556_),
    .A2(_2498_),
    .ZN(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7303_ (.A1(_2498_),
    .A2(_2502_),
    .B(_2503_),
    .C(_2127_),
    .ZN(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7304_ (.A1(_0454_),
    .A2(_0475_),
    .Z(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7305_ (.A1(_2450_),
    .A2(_2451_),
    .B(_2505_),
    .ZN(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7306_ (.A1(_0556_),
    .A2(_0575_),
    .A3(_2506_),
    .Z(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7307_ (.A1(_1555_),
    .A2(_2358_),
    .ZN(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7308_ (.A1(_2358_),
    .A2(_2507_),
    .B(_2508_),
    .C(_2135_),
    .ZN(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7309_ (.A1(_2350_),
    .A2(_2504_),
    .A3(_2509_),
    .ZN(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7310_ (.A1(_2497_),
    .A2(_2510_),
    .ZN(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7311_ (.A1(_2491_),
    .A2(net9),
    .ZN(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7312_ (.A1(_2491_),
    .A2(net9),
    .Z(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7313_ (.A1(_2512_),
    .A2(_2513_),
    .ZN(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7314_ (.A1(_1073_),
    .A2(_0453_),
    .ZN(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7315_ (.A1(_2515_),
    .A2(_2462_),
    .Z(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7316_ (.A1(_2514_),
    .A2(_2516_),
    .ZN(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7317_ (.A1(_2496_),
    .A2(_2511_),
    .B1(_2517_),
    .B2(_2153_),
    .ZN(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7318_ (.A1(_1084_),
    .A2(_2419_),
    .ZN(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7319_ (.A1(_2459_),
    .A2(_2481_),
    .ZN(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7320_ (.A1(_2515_),
    .A2(_2520_),
    .ZN(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7321_ (.A1(_2514_),
    .A2(_2521_),
    .Z(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7322_ (.I(net53),
    .ZN(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7323_ (.A1(_2523_),
    .A2(_2323_),
    .ZN(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7324_ (.A1(_1545_),
    .A2(_2522_),
    .B(_2524_),
    .C(_2421_),
    .ZN(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7325_ (.I(_0936_),
    .Z(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7326_ (.I(_2474_),
    .Z(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7327_ (.I(_2340_),
    .Z(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7328_ (.A1(_2528_),
    .A2(_2495_),
    .B(_2345_),
    .ZN(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7329_ (.A1(net53),
    .A2(_2526_),
    .B1(_2527_),
    .B2(_1556_),
    .C(_2529_),
    .ZN(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7330_ (.I(_1155_),
    .Z(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7331_ (.A1(_2525_),
    .A2(_2530_),
    .B(_2531_),
    .ZN(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7332_ (.I(_1676_),
    .Z(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7333_ (.A1(_2519_),
    .A2(_2532_),
    .B(_2533_),
    .ZN(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7334_ (.A1(_1084_),
    .A2(_2239_),
    .B1(_1488_),
    .B2(_2518_),
    .C(_2534_),
    .ZN(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7335_ (.I(_2382_),
    .Z(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7336_ (.A1(_2492_),
    .A2(_2493_),
    .B1(_2535_),
    .B2(_2536_),
    .ZN(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7337_ (.A1(net53),
    .A2(_2377_),
    .B(_1425_),
    .ZN(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7338_ (.A1(_2307_),
    .A2(_2537_),
    .B(_2538_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7339_ (.I(\as2650.pc[4] ),
    .Z(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7340_ (.I(_2539_),
    .Z(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7341_ (.I(_2540_),
    .Z(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7342_ (.I(_2350_),
    .Z(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7343_ (.I(_0554_),
    .Z(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7344_ (.A1(_2543_),
    .A2(_1271_),
    .ZN(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7345_ (.A1(_2543_),
    .A2(_1271_),
    .B1(_2443_),
    .B2(_2499_),
    .C(_2500_),
    .ZN(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7346_ (.A1(_2544_),
    .A2(_2545_),
    .ZN(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7347_ (.A1(_1288_),
    .A2(_0643_),
    .A3(_2546_),
    .ZN(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7348_ (.A1(_2387_),
    .A2(_2547_),
    .ZN(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7349_ (.A1(_1558_),
    .A2(_2387_),
    .B(_2354_),
    .C(_2548_),
    .ZN(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7350_ (.A1(_2543_),
    .A2(_0574_),
    .ZN(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7351_ (.A1(_2543_),
    .A2(_0574_),
    .B1(_2450_),
    .B2(_2451_),
    .C(_2505_),
    .ZN(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7352_ (.A1(_2550_),
    .A2(_2551_),
    .ZN(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7353_ (.A1(_1288_),
    .A2(_0686_),
    .A3(_2552_),
    .ZN(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7354_ (.A1(_2395_),
    .A2(_2553_),
    .ZN(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7355_ (.A1(_1558_),
    .A2(_2395_),
    .B(_2554_),
    .C(_2399_),
    .ZN(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7356_ (.A1(_2549_),
    .A2(_2555_),
    .ZN(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7357_ (.I(_1487_),
    .Z(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7358_ (.A1(_2539_),
    .A2(_0674_),
    .Z(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7359_ (.A1(_2492_),
    .A2(_0555_),
    .ZN(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7360_ (.A1(_2512_),
    .A2(_2516_),
    .B(_2559_),
    .ZN(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7361_ (.A1(_2558_),
    .A2(_2560_),
    .ZN(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _7362_ (.I(_2366_),
    .ZN(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7363_ (.A1(_2562_),
    .A2(_2351_),
    .ZN(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7364_ (.A1(_2558_),
    .A2(_2560_),
    .ZN(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7365_ (.A1(_2563_),
    .A2(_2564_),
    .ZN(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7366_ (.I(net32),
    .Z(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7367_ (.A1(_2523_),
    .A2(_2494_),
    .ZN(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7368_ (.A1(_2566_),
    .A2(_2567_),
    .Z(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7369_ (.A1(_2561_),
    .A2(_2565_),
    .B1(_2568_),
    .B2(_2466_),
    .ZN(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7370_ (.A1(_2557_),
    .A2(_2569_),
    .ZN(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7371_ (.A1(_2542_),
    .A2(_2556_),
    .B(_2570_),
    .ZN(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7372_ (.A1(_2209_),
    .A2(_1415_),
    .ZN(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7373_ (.I(_2572_),
    .Z(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7374_ (.I(_2417_),
    .Z(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7375_ (.A1(_2573_),
    .A2(_2574_),
    .ZN(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7376_ (.A1(_2566_),
    .A2(_2472_),
    .B(_2346_),
    .ZN(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7377_ (.I(_2413_),
    .Z(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7378_ (.I(_2475_),
    .Z(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7379_ (.A1(_1558_),
    .A2(_2577_),
    .B1(_2568_),
    .B2(_2578_),
    .ZN(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7380_ (.I(_2512_),
    .ZN(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _7381_ (.A1(_2580_),
    .A2(_2521_),
    .B(_2513_),
    .ZN(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7382_ (.A1(_2558_),
    .A2(_2581_),
    .Z(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7383_ (.A1(_2321_),
    .A2(_2582_),
    .ZN(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7384_ (.A1(_2566_),
    .A2(_2324_),
    .B(_2329_),
    .C(_2583_),
    .ZN(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7385_ (.A1(_2576_),
    .A2(_2579_),
    .B(_2584_),
    .ZN(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7386_ (.I(_2573_),
    .Z(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7387_ (.I(_1631_),
    .Z(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7388_ (.I(_2587_),
    .Z(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7389_ (.A1(_2541_),
    .A2(_2575_),
    .B1(_2585_),
    .B2(_2586_),
    .C(_2588_),
    .ZN(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7390_ (.A1(_2571_),
    .A2(_2589_),
    .B(_2374_),
    .ZN(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7391_ (.A1(_2541_),
    .A2(_2493_),
    .B(_2590_),
    .ZN(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7392_ (.A1(_2566_),
    .A2(_2377_),
    .B(_1425_),
    .ZN(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7393_ (.A1(_2307_),
    .A2(_2591_),
    .B(_2592_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7394_ (.I(\as2650.pc[5] ),
    .Z(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7395_ (.I(_2593_),
    .Z(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7396_ (.I(_2594_),
    .Z(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7397_ (.I(_4256_),
    .Z(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7398_ (.A1(net32),
    .A2(_2567_),
    .Z(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7399_ (.A1(net33),
    .A2(_2597_),
    .Z(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7400_ (.A1(_2596_),
    .A2(_2598_),
    .ZN(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7401_ (.I(net33),
    .Z(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7402_ (.I(_2136_),
    .Z(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7403_ (.A1(_2600_),
    .A2(_0936_),
    .B(_2344_),
    .C(_2601_),
    .ZN(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7404_ (.A1(_2179_),
    .A2(_2413_),
    .B(_2599_),
    .C(_2602_),
    .ZN(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7405_ (.I(_1581_),
    .Z(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7406_ (.I(_2604_),
    .Z(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7407_ (.I(net1),
    .Z(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7408_ (.A1(_2593_),
    .A2(_2606_),
    .Z(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7409_ (.A1(_1091_),
    .A2(net10),
    .Z(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7410_ (.A1(_2608_),
    .A2(_2581_),
    .ZN(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7411_ (.A1(_2540_),
    .A2(_0675_),
    .B(_2609_),
    .ZN(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7412_ (.A1(_2607_),
    .A2(_2610_),
    .Z(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7413_ (.A1(_2600_),
    .A2(_2185_),
    .ZN(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7414_ (.A1(_2605_),
    .A2(_2611_),
    .B(_2612_),
    .C(_2328_),
    .ZN(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7415_ (.A1(_2603_),
    .A2(_2613_),
    .ZN(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7416_ (.I(_1189_),
    .Z(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7417_ (.A1(_1097_),
    .A2(_2419_),
    .B1(_2614_),
    .B2(_2615_),
    .ZN(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7418_ (.A1(_2366_),
    .A2(_2152_),
    .Z(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7419_ (.A1(_1096_),
    .A2(_0755_),
    .Z(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7420_ (.A1(_2539_),
    .A2(net10),
    .ZN(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7421_ (.A1(_2619_),
    .A2(_2561_),
    .ZN(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7422_ (.A1(_2618_),
    .A2(_2620_),
    .Z(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7423_ (.A1(_2606_),
    .A2(_0740_),
    .Z(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7424_ (.I(net10),
    .Z(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7425_ (.A1(_2623_),
    .A2(_0685_),
    .ZN(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7426_ (.A1(_2623_),
    .A2(_0685_),
    .ZN(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _7427_ (.A1(_2550_),
    .A2(_2624_),
    .A3(_2551_),
    .B(_2625_),
    .ZN(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7428_ (.A1(_2622_),
    .A2(_2626_),
    .Z(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7429_ (.A1(_2622_),
    .A2(_2626_),
    .B(_2357_),
    .ZN(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7430_ (.I(_4242_),
    .Z(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7431_ (.A1(_1410_),
    .A2(_2357_),
    .B1(_2627_),
    .B2(_2628_),
    .C(_2629_),
    .ZN(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7432_ (.A1(_2623_),
    .A2(_0642_),
    .ZN(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7433_ (.A1(_2623_),
    .A2(_0642_),
    .ZN(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _7434_ (.A1(_2544_),
    .A2(_2631_),
    .A3(_2545_),
    .B(_2632_),
    .ZN(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7435_ (.A1(_0757_),
    .A2(_0771_),
    .A3(_2633_),
    .Z(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7436_ (.A1(_1585_),
    .A2(_4447_),
    .B(_2126_),
    .ZN(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7437_ (.A1(_2389_),
    .A2(_2634_),
    .B(_2635_),
    .ZN(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7438_ (.A1(_2351_),
    .A2(_2630_),
    .A3(_2636_),
    .B(_2497_),
    .ZN(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7439_ (.A1(_2402_),
    .A2(_2598_),
    .B(_2637_),
    .ZN(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7440_ (.A1(_2617_),
    .A2(_2621_),
    .B(_2638_),
    .C(_2439_),
    .ZN(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7441_ (.A1(_2595_),
    .A2(_2438_),
    .B1(_2533_),
    .B2(_2616_),
    .C(_2639_),
    .ZN(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7442_ (.A1(_2309_),
    .A2(_2640_),
    .ZN(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7443_ (.A1(_2595_),
    .A2(_2493_),
    .B(_2641_),
    .ZN(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7444_ (.I(_2305_),
    .Z(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7445_ (.I(_1424_),
    .Z(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7446_ (.A1(_2600_),
    .A2(_2643_),
    .B(_2644_),
    .ZN(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7447_ (.A1(_2307_),
    .A2(_2642_),
    .B(_2645_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7448_ (.I(_2434_),
    .Z(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7449_ (.I(_1103_),
    .Z(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7450_ (.I(_2629_),
    .Z(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7451_ (.I(_0830_),
    .Z(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7452_ (.A1(_2649_),
    .A2(_0840_),
    .ZN(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7453_ (.A1(_0756_),
    .A2(_0741_),
    .Z(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7454_ (.A1(_2622_),
    .A2(_2626_),
    .B(_2651_),
    .ZN(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7455_ (.A1(_2650_),
    .A2(_2652_),
    .B(_2394_),
    .ZN(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7456_ (.A1(_2650_),
    .A2(_2652_),
    .B(_2653_),
    .ZN(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7457_ (.A1(_1560_),
    .A2(_2358_),
    .B(_2654_),
    .ZN(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7458_ (.A1(_1596_),
    .A2(_0820_),
    .ZN(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7459_ (.A1(_0756_),
    .A2(_0770_),
    .Z(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7460_ (.A1(_0756_),
    .A2(_0770_),
    .Z(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7461_ (.A1(_2633_),
    .A2(_2657_),
    .B(_2658_),
    .ZN(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7462_ (.A1(_2656_),
    .A2(_2659_),
    .ZN(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7463_ (.A1(_2389_),
    .A2(_2660_),
    .ZN(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7464_ (.A1(_1559_),
    .A2(_2387_),
    .B(_2354_),
    .C(_2661_),
    .ZN(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7465_ (.A1(_2648_),
    .A2(_2655_),
    .B(_2662_),
    .ZN(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7466_ (.A1(_2558_),
    .A2(_2560_),
    .A3(_2607_),
    .ZN(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7467_ (.A1(_1096_),
    .A2(_1584_),
    .B(_2619_),
    .ZN(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7468_ (.A1(_2593_),
    .A2(_0755_),
    .B(_2665_),
    .ZN(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7469_ (.A1(_1105_),
    .A2(_1597_),
    .Z(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7470_ (.A1(_2664_),
    .A2(_2666_),
    .B(_2667_),
    .ZN(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7471_ (.A1(_2667_),
    .A2(_2664_),
    .A3(_2666_),
    .ZN(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7472_ (.A1(_2368_),
    .A2(_2669_),
    .ZN(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7473_ (.I(net34),
    .Z(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7474_ (.A1(_2600_),
    .A2(_2597_),
    .ZN(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7475_ (.A1(_2671_),
    .A2(_2672_),
    .ZN(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7476_ (.A1(_2466_),
    .A2(_2673_),
    .ZN(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7477_ (.A1(_2668_),
    .A2(_2670_),
    .B(_2674_),
    .ZN(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7478_ (.A1(_2542_),
    .A2(_2663_),
    .B(_2675_),
    .C(_2386_),
    .ZN(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7479_ (.I(_2236_),
    .Z(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7480_ (.A1(_2677_),
    .A2(_2673_),
    .ZN(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7481_ (.A1(_2671_),
    .A2(_2472_),
    .B1(_2577_),
    .B2(_1559_),
    .C(_2346_),
    .ZN(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7482_ (.A1(_2608_),
    .A2(_2581_),
    .A3(_2618_),
    .B(_2666_),
    .ZN(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7483_ (.A1(_2667_),
    .A2(_2680_),
    .Z(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7484_ (.A1(_2321_),
    .A2(_2681_),
    .ZN(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7485_ (.A1(_2671_),
    .A2(_2324_),
    .B(_2329_),
    .C(_2682_),
    .ZN(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7486_ (.A1(_2678_),
    .A2(_2679_),
    .B(_2683_),
    .ZN(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7487_ (.A1(_2647_),
    .A2(_2575_),
    .B1(_2684_),
    .B2(_2586_),
    .C(_2588_),
    .ZN(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7488_ (.A1(_2676_),
    .A2(_2685_),
    .B(_2374_),
    .ZN(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7489_ (.A1(_2647_),
    .A2(_2493_),
    .B(_2686_),
    .ZN(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7490_ (.A1(_2671_),
    .A2(_2643_),
    .B(_2644_),
    .ZN(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7491_ (.A1(_2646_),
    .A2(_2687_),
    .B(_2688_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7492_ (.I(_1110_),
    .Z(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7493_ (.I(net35),
    .Z(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7494_ (.A1(net34),
    .A2(net33),
    .A3(_2597_),
    .ZN(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7495_ (.A1(_2690_),
    .A2(_2691_),
    .Z(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7496_ (.A1(_2690_),
    .A2(_2526_),
    .B1(_2474_),
    .B2(_2321_),
    .ZN(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7497_ (.A1(_1658_),
    .A2(_0940_),
    .ZN(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7498_ (.I(_2694_),
    .Z(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7499_ (.A1(_2578_),
    .A2(_2692_),
    .B(_2693_),
    .C(_2695_),
    .ZN(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7500_ (.A1(_2689_),
    .A2(_2316_),
    .B(_2696_),
    .ZN(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7501_ (.A1(\as2650.pc[7] ),
    .A2(net2),
    .Z(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7502_ (.A1(_1103_),
    .A2(_1595_),
    .ZN(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7503_ (.A1(\as2650.pc[6] ),
    .A2(net2),
    .Z(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7504_ (.A1(_2700_),
    .A2(_2680_),
    .ZN(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7505_ (.A1(_2699_),
    .A2(_2701_),
    .ZN(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7506_ (.A1(_2698_),
    .A2(_2702_),
    .Z(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7507_ (.A1(_2690_),
    .A2(_2605_),
    .ZN(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7508_ (.A1(_2222_),
    .A2(_1572_),
    .A3(_2423_),
    .A4(_2704_),
    .ZN(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7509_ (.A1(_2322_),
    .A2(_2703_),
    .B(_2705_),
    .ZN(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7510_ (.A1(_2647_),
    .A2(_1525_),
    .B(_2668_),
    .ZN(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7511_ (.A1(_2698_),
    .A2(_2707_),
    .ZN(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7512_ (.A1(_1597_),
    .A2(_0841_),
    .ZN(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7513_ (.A1(_2650_),
    .A2(_2652_),
    .B(_2709_),
    .ZN(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7514_ (.A1(_1599_),
    .A2(_0893_),
    .A3(_2710_),
    .Z(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7515_ (.A1(_4428_),
    .A2(_2711_),
    .ZN(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7516_ (.A1(_2185_),
    .A2(_2394_),
    .B(_2712_),
    .C(_2134_),
    .ZN(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7517_ (.A1(_0831_),
    .A2(_0821_),
    .ZN(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7518_ (.A1(_2656_),
    .A2(_2659_),
    .B(_2714_),
    .ZN(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7519_ (.A1(_0933_),
    .A2(_0891_),
    .A3(_2715_),
    .Z(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7520_ (.A1(_2320_),
    .A2(_2498_),
    .ZN(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7521_ (.A1(_2498_),
    .A2(_2716_),
    .B(_2717_),
    .C(_2353_),
    .ZN(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7522_ (.I(_2497_),
    .ZN(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7523_ (.A1(_2713_),
    .A2(_2718_),
    .B(_2719_),
    .ZN(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7524_ (.A1(_2466_),
    .A2(_2692_),
    .B(_2720_),
    .C(_2405_),
    .ZN(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7525_ (.A1(_2153_),
    .A2(_2708_),
    .B(_2721_),
    .C(_2385_),
    .ZN(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7526_ (.A1(_2317_),
    .A2(_2697_),
    .B(_2706_),
    .C(_2722_),
    .ZN(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7527_ (.I(_2382_),
    .Z(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7528_ (.A1(_2689_),
    .A2(_2384_),
    .B1(_2723_),
    .B2(_2724_),
    .ZN(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7529_ (.A1(_2690_),
    .A2(_2434_),
    .ZN(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7530_ (.A1(_2377_),
    .A2(_2725_),
    .B(_2726_),
    .C(_2437_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7531_ (.I(_2383_),
    .Z(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7532_ (.A1(_1599_),
    .A2(_0893_),
    .ZN(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7533_ (.A1(_2650_),
    .A2(_2652_),
    .B(_2728_),
    .C(_2709_),
    .ZN(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7534_ (.I(_2729_),
    .Z(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7535_ (.A1(_1336_),
    .A2(_0894_),
    .Z(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7536_ (.A1(_4428_),
    .A2(_2731_),
    .Z(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7537_ (.A1(_2730_),
    .A2(_2732_),
    .ZN(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7538_ (.A1(_2161_),
    .A2(_2733_),
    .Z(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7539_ (.I(_2160_),
    .ZN(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7540_ (.A1(_0900_),
    .A2(_0890_),
    .ZN(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7541_ (.A1(_2656_),
    .A2(_2659_),
    .B(_2736_),
    .C(_2714_),
    .ZN(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7542_ (.A1(_1599_),
    .A2(_0890_),
    .ZN(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7543_ (.A1(_4277_),
    .A2(_2738_),
    .ZN(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7544_ (.A1(_2737_),
    .A2(_2739_),
    .Z(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7545_ (.I(_2740_),
    .Z(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7546_ (.A1(_2735_),
    .A2(_2741_),
    .Z(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7547_ (.A1(_2362_),
    .A2(_2734_),
    .B1(_2742_),
    .B2(_2354_),
    .ZN(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7548_ (.I(net36),
    .Z(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7549_ (.I(net35),
    .ZN(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7550_ (.A1(_2745_),
    .A2(_2691_),
    .ZN(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7551_ (.A1(_2744_),
    .A2(_2746_),
    .ZN(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7552_ (.I(_2405_),
    .Z(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7553_ (.A1(_2365_),
    .A2(_2747_),
    .B(_2748_),
    .ZN(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7554_ (.A1(_2352_),
    .A2(_2743_),
    .B(_2749_),
    .ZN(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7555_ (.A1(\as2650.pc[8] ),
    .A2(_1595_),
    .Z(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7556_ (.A1(_2700_),
    .A2(_2698_),
    .ZN(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7557_ (.A1(_1110_),
    .A2(_0830_),
    .ZN(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7558_ (.A1(_2666_),
    .A2(_2752_),
    .B(_2753_),
    .C(_2699_),
    .ZN(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7559_ (.A1(_2664_),
    .A2(_2752_),
    .ZN(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7560_ (.A1(_2754_),
    .A2(_2755_),
    .Z(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7561_ (.A1(_2751_),
    .A2(_2756_),
    .ZN(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7562_ (.I(_2563_),
    .Z(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7563_ (.A1(_2751_),
    .A2(_2756_),
    .ZN(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7564_ (.A1(_2758_),
    .A2(_2759_),
    .ZN(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7565_ (.A1(_2757_),
    .A2(_2760_),
    .B(_2386_),
    .ZN(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7566_ (.A1(_2744_),
    .A2(_2341_),
    .B1(_2577_),
    .B2(_2162_),
    .C(_2345_),
    .ZN(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7567_ (.A1(_0409_),
    .A2(_2747_),
    .B(_2762_),
    .ZN(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _7568_ (.A1(_2608_),
    .A2(_2581_),
    .A3(_2618_),
    .A4(_2752_),
    .ZN(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7569_ (.A1(_2754_),
    .A2(_2764_),
    .B(_2751_),
    .ZN(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _7570_ (.A1(_2751_),
    .A2(_2754_),
    .A3(_2764_),
    .Z(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7571_ (.A1(_2765_),
    .A2(_2766_),
    .ZN(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7572_ (.I(_2426_),
    .Z(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7573_ (.A1(_2744_),
    .A2(_2768_),
    .ZN(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7574_ (.A1(_2322_),
    .A2(_2767_),
    .B(_2769_),
    .C(_2421_),
    .ZN(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7575_ (.A1(_2763_),
    .A2(_2770_),
    .B(_2586_),
    .ZN(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7576_ (.I(_1631_),
    .Z(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7577_ (.A1(_0968_),
    .A2(_2575_),
    .B(_2772_),
    .ZN(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7578_ (.A1(_2750_),
    .A2(_2761_),
    .B1(_2771_),
    .B2(_2773_),
    .ZN(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7579_ (.A1(_0968_),
    .A2(_2727_),
    .B1(_2774_),
    .B2(_2536_),
    .ZN(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7580_ (.A1(_2744_),
    .A2(_2643_),
    .B(_2644_),
    .ZN(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7581_ (.A1(_2646_),
    .A2(_2775_),
    .B(_2776_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7582_ (.I(\as2650.pc[9] ),
    .Z(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7583_ (.I(_2334_),
    .Z(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7584_ (.I(_2778_),
    .Z(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7585_ (.I(net37),
    .Z(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7586_ (.A1(net36),
    .A2(_2746_),
    .ZN(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7587_ (.A1(_2780_),
    .A2(_2781_),
    .Z(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7588_ (.A1(_2779_),
    .A2(_2782_),
    .ZN(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7589_ (.A1(_2165_),
    .A2(_2778_),
    .ZN(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7590_ (.A1(_2780_),
    .A2(_2526_),
    .ZN(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7591_ (.A1(_2332_),
    .A2(_2784_),
    .B(_2785_),
    .C(_2695_),
    .ZN(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7592_ (.A1(_2777_),
    .A2(_2316_),
    .B1(_2783_),
    .B2(_2786_),
    .ZN(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7593_ (.A1(_0985_),
    .A2(_1595_),
    .Z(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7594_ (.I(_2788_),
    .Z(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7595_ (.A1(_0966_),
    .A2(_0832_),
    .ZN(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7596_ (.A1(_2790_),
    .A2(_2765_),
    .ZN(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7597_ (.A1(_2789_),
    .A2(_2791_),
    .ZN(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7598_ (.I(_2185_),
    .Z(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7599_ (.A1(_2780_),
    .A2(_2793_),
    .Z(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7600_ (.A1(_1420_),
    .A2(_2329_),
    .ZN(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7601_ (.A1(_1691_),
    .A2(_2792_),
    .B(_2794_),
    .C(_2795_),
    .ZN(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7602_ (.I(_1477_),
    .Z(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7603_ (.A1(_2161_),
    .A2(_2165_),
    .A3(_2741_),
    .ZN(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7604_ (.A1(_2388_),
    .A2(_2798_),
    .ZN(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7605_ (.A1(_2162_),
    .A2(_2741_),
    .B(_2165_),
    .ZN(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7606_ (.A1(_2160_),
    .A2(\as2650.addr_buff[1] ),
    .A3(_2730_),
    .A4(_2732_),
    .Z(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7607_ (.A1(_2629_),
    .A2(_2801_),
    .ZN(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _7608_ (.I(\as2650.addr_buff[1] ),
    .ZN(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7609_ (.A1(_2735_),
    .A2(_2733_),
    .B(_2803_),
    .ZN(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7610_ (.A1(_2802_),
    .A2(_2804_),
    .ZN(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7611_ (.A1(_2799_),
    .A2(_2800_),
    .B(_2805_),
    .ZN(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7612_ (.A1(_2790_),
    .A2(_2757_),
    .ZN(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7613_ (.A1(_2789_),
    .A2(_2807_),
    .Z(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7614_ (.A1(_2758_),
    .A2(_2808_),
    .B1(_2782_),
    .B2(_2402_),
    .ZN(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7615_ (.A1(_2542_),
    .A2(_2806_),
    .B(_2809_),
    .C(_2385_),
    .ZN(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7616_ (.A1(_1573_),
    .A2(_2787_),
    .B1(_2796_),
    .B2(_2797_),
    .C(_2810_),
    .ZN(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7617_ (.A1(_2777_),
    .A2(_2727_),
    .B1(_2811_),
    .B2(_2536_),
    .ZN(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7618_ (.A1(_2780_),
    .A2(_2643_),
    .B(_2644_),
    .ZN(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7619_ (.A1(_2646_),
    .A2(_2812_),
    .B(_2813_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7620_ (.I(\as2650.pc[10] ),
    .Z(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7621_ (.I(_2814_),
    .Z(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7622_ (.I(net52),
    .ZN(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7623_ (.A1(net37),
    .A2(net36),
    .A3(_2746_),
    .ZN(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7624_ (.A1(_2816_),
    .A2(_2817_),
    .Z(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7625_ (.A1(_2388_),
    .A2(_2798_),
    .B(_2802_),
    .ZN(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7626_ (.A1(\as2650.addr_buff[0] ),
    .A2(\as2650.addr_buff[1] ),
    .A3(\as2650.addr_buff[2] ),
    .Z(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7627_ (.I(_2820_),
    .Z(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7628_ (.A1(_4248_),
    .A2(_2731_),
    .A3(_2730_),
    .ZN(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7629_ (.A1(_2353_),
    .A2(_2737_),
    .A3(_2739_),
    .ZN(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7630_ (.A1(_2822_),
    .A2(_2823_),
    .ZN(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7631_ (.A1(_2821_),
    .A2(_2824_),
    .ZN(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7632_ (.A1(_2169_),
    .A2(_2819_),
    .B(_2825_),
    .ZN(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7633_ (.A1(_2542_),
    .A2(_2826_),
    .ZN(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7634_ (.A1(_2402_),
    .A2(_2818_),
    .B(_2827_),
    .C(_2758_),
    .ZN(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7635_ (.A1(_0997_),
    .A2(_0830_),
    .Z(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7636_ (.I(_2829_),
    .Z(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7637_ (.A1(_2777_),
    .A2(\as2650.pc[8] ),
    .B(_2649_),
    .ZN(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7638_ (.I(_2831_),
    .ZN(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7639_ (.A1(_2757_),
    .A2(_2789_),
    .ZN(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7640_ (.A1(_2832_),
    .A2(_2833_),
    .ZN(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7641_ (.A1(_2830_),
    .A2(_2834_),
    .Z(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7642_ (.A1(_2153_),
    .A2(_2835_),
    .B(_2386_),
    .ZN(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7643_ (.A1(_1475_),
    .A2(_1663_),
    .ZN(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7644_ (.I(_2837_),
    .Z(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7645_ (.I(_2838_),
    .Z(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7646_ (.A1(_2677_),
    .A2(_2818_),
    .ZN(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7647_ (.I(_1443_),
    .Z(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7648_ (.A1(net52),
    .A2(_2472_),
    .B1(_2577_),
    .B2(_2169_),
    .C(_2841_),
    .ZN(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7649_ (.A1(_0998_),
    .A2(_2574_),
    .B1(_2840_),
    .B2(_2842_),
    .ZN(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7650_ (.A1(_2839_),
    .A2(_2843_),
    .ZN(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7651_ (.A1(_2765_),
    .A2(_2788_),
    .B(_2831_),
    .ZN(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7652_ (.A1(_2830_),
    .A2(_2845_),
    .Z(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7653_ (.A1(net52),
    .A2(_2768_),
    .B(_2423_),
    .ZN(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7654_ (.A1(_2322_),
    .A2(_2846_),
    .B(_2847_),
    .ZN(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7655_ (.A1(_2815_),
    .A2(_2348_),
    .B1(_2848_),
    .B2(_2223_),
    .C(_2772_),
    .ZN(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7656_ (.A1(_2828_),
    .A2(_2836_),
    .B1(_2844_),
    .B2(_2849_),
    .ZN(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7657_ (.A1(_2815_),
    .A2(_2727_),
    .B1(_2850_),
    .B2(_2536_),
    .ZN(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7658_ (.I(_1424_),
    .Z(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7659_ (.A1(net52),
    .A2(_2306_),
    .B(_2852_),
    .ZN(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7660_ (.A1(_2646_),
    .A2(_2851_),
    .B(_2853_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7661_ (.I(\as2650.pc[11] ),
    .Z(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7662_ (.I(_2854_),
    .Z(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7663_ (.I(_2855_),
    .Z(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7664_ (.I(net39),
    .Z(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7665_ (.A1(_2816_),
    .A2(_2817_),
    .ZN(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7666_ (.A1(_2857_),
    .A2(_2858_),
    .ZN(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7667_ (.A1(_2730_),
    .A2(_2732_),
    .A3(_2821_),
    .ZN(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7668_ (.A1(_2741_),
    .A2(_2821_),
    .ZN(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7669_ (.A1(_2135_),
    .A2(_2860_),
    .B1(_2861_),
    .B2(_2127_),
    .C(_2172_),
    .ZN(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7670_ (.A1(_2173_),
    .A2(_2825_),
    .B(_2862_),
    .C(_2719_),
    .ZN(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7671_ (.A1(_2365_),
    .A2(_2859_),
    .B(_2863_),
    .C(_2368_),
    .ZN(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7672_ (.A1(_1008_),
    .A2(_1596_),
    .Z(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7673_ (.A1(_2814_),
    .A2(_2649_),
    .ZN(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7674_ (.A1(_2830_),
    .A2(_2834_),
    .B(_2866_),
    .ZN(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7675_ (.A1(_2865_),
    .A2(_2867_),
    .Z(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7676_ (.A1(_2617_),
    .A2(_2868_),
    .ZN(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7677_ (.A1(_2864_),
    .A2(_2869_),
    .ZN(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7678_ (.A1(_2857_),
    .A2(_2526_),
    .B1(_2527_),
    .B2(_2173_),
    .ZN(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7679_ (.A1(_2578_),
    .A2(_2859_),
    .B(_2871_),
    .C(_2695_),
    .ZN(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7680_ (.I(_2312_),
    .Z(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7681_ (.A1(_2856_),
    .A2(_2574_),
    .ZN(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7682_ (.A1(_1008_),
    .A2(_2873_),
    .B1(_2874_),
    .B2(_2838_),
    .ZN(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7683_ (.A1(_2872_),
    .A2(_2875_),
    .B(_2772_),
    .ZN(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7684_ (.I(_2845_),
    .ZN(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7685_ (.A1(_2830_),
    .A2(_2877_),
    .B(_2866_),
    .ZN(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7686_ (.A1(_2865_),
    .A2(_2878_),
    .ZN(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7687_ (.A1(_2768_),
    .A2(_2879_),
    .ZN(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7688_ (.A1(_2423_),
    .A2(_2880_),
    .ZN(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7689_ (.A1(_2857_),
    .A2(_2186_),
    .B(_1676_),
    .C(_2881_),
    .ZN(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7690_ (.A1(_1488_),
    .A2(_2870_),
    .B(_2876_),
    .C(_2882_),
    .ZN(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7691_ (.A1(_2856_),
    .A2(_2727_),
    .B1(_2883_),
    .B2(_2724_),
    .ZN(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7692_ (.A1(_2857_),
    .A2(_2306_),
    .B(_2852_),
    .ZN(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7693_ (.A1(_2379_),
    .A2(_2884_),
    .B(_2885_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7694_ (.I(\as2650.pc[12] ),
    .Z(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7695_ (.A1(_2829_),
    .A2(_2865_),
    .ZN(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7696_ (.A1(\as2650.pc[11] ),
    .A2(_0831_),
    .ZN(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7697_ (.A1(_2866_),
    .A2(_2831_),
    .A3(_2888_),
    .ZN(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7698_ (.A1(_2833_),
    .A2(_2887_),
    .B(_2889_),
    .ZN(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7699_ (.A1(\as2650.pc[12] ),
    .A2(_0831_),
    .Z(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7700_ (.A1(_2890_),
    .A2(_2891_),
    .Z(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7701_ (.A1(\as2650.addr_buff[3] ),
    .A2(_2729_),
    .A3(_2732_),
    .A4(_2820_),
    .ZN(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7702_ (.A1(_2177_),
    .A2(_2893_),
    .Z(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7703_ (.A1(\as2650.addr_buff[3] ),
    .A2(_2740_),
    .A3(_2821_),
    .ZN(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7704_ (.A1(_2177_),
    .A2(_2895_),
    .Z(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7705_ (.A1(_2361_),
    .A2(_2894_),
    .B1(_2896_),
    .B2(_2388_),
    .ZN(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7706_ (.A1(net39),
    .A2(_2858_),
    .ZN(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7707_ (.A1(net51),
    .A2(_2898_),
    .Z(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7708_ (.A1(_2364_),
    .A2(_2899_),
    .ZN(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7709_ (.A1(_2352_),
    .A2(_2897_),
    .B(_2900_),
    .C(_2758_),
    .ZN(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7710_ (.A1(_2617_),
    .A2(_2892_),
    .B(_2901_),
    .C(_2370_),
    .ZN(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7711_ (.I(\as2650.addr_buff[4] ),
    .ZN(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7712_ (.A1(_2903_),
    .A2(_2338_),
    .ZN(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7713_ (.A1(net51),
    .A2(_0936_),
    .B1(_2904_),
    .B2(_2187_),
    .ZN(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7714_ (.A1(_2476_),
    .A2(_2899_),
    .B(_2905_),
    .C(_2695_),
    .ZN(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7715_ (.A1(_2886_),
    .A2(_2316_),
    .B(_2906_),
    .ZN(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7716_ (.A1(_2765_),
    .A2(_2789_),
    .ZN(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7717_ (.A1(_2908_),
    .A2(_2887_),
    .B(_2889_),
    .ZN(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7718_ (.A1(_2891_),
    .A2(_2909_),
    .Z(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7719_ (.A1(_2793_),
    .A2(_2910_),
    .ZN(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7720_ (.A1(net51),
    .A2(_2793_),
    .B(_2795_),
    .C(_2911_),
    .ZN(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7721_ (.A1(_1513_),
    .A2(_2907_),
    .B1(_2912_),
    .B2(_1477_),
    .ZN(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7722_ (.A1(_2902_),
    .A2(_2913_),
    .Z(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7723_ (.A1(_2886_),
    .A2(_2384_),
    .B1(_2914_),
    .B2(_2724_),
    .ZN(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7724_ (.A1(net51),
    .A2(_2306_),
    .B(_2852_),
    .ZN(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7725_ (.A1(_2379_),
    .A2(_2915_),
    .B(_2916_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7726_ (.A1(_1324_),
    .A2(_2381_),
    .ZN(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7727_ (.A1(_2320_),
    .A2(_2367_),
    .ZN(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7728_ (.I(_2918_),
    .ZN(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7729_ (.A1(_1486_),
    .A2(_2125_),
    .B1(_2917_),
    .B2(_2919_),
    .ZN(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7730_ (.A1(_1387_),
    .A2(_2273_),
    .B(_1473_),
    .ZN(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7731_ (.A1(_4427_),
    .A2(_4425_),
    .ZN(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7732_ (.A1(_4420_),
    .A2(_2922_),
    .ZN(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7733_ (.A1(_1466_),
    .A2(_4170_),
    .B(_2923_),
    .ZN(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7734_ (.A1(_2238_),
    .A2(_2920_),
    .A3(_2921_),
    .A4(_2924_),
    .ZN(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7735_ (.A1(_1032_),
    .A2(_1375_),
    .A3(_2257_),
    .Z(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7736_ (.A1(_2281_),
    .A2(_2284_),
    .ZN(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7737_ (.A1(_2243_),
    .A2(_2927_),
    .A3(_2292_),
    .ZN(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7738_ (.A1(_1657_),
    .A2(_1664_),
    .B1(_2917_),
    .B2(_2719_),
    .C(_2928_),
    .ZN(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7739_ (.A1(_2255_),
    .A2(_2262_),
    .A3(_2926_),
    .A4(_2929_),
    .ZN(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7740_ (.A1(_2268_),
    .A2(_2925_),
    .A3(_2930_),
    .ZN(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7741_ (.A1(_2290_),
    .A2(_2931_),
    .ZN(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7742_ (.A1(_2303_),
    .A2(_2932_),
    .ZN(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7743_ (.I(_2150_),
    .Z(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7744_ (.I(_2934_),
    .Z(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7745_ (.A1(net50),
    .A2(_2615_),
    .ZN(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7746_ (.A1(_2935_),
    .A2(_2936_),
    .ZN(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7747_ (.A1(_1574_),
    .A2(_2936_),
    .B(_2203_),
    .C(_2239_),
    .ZN(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7748_ (.I(_2244_),
    .Z(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7749_ (.I(_2939_),
    .Z(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7750_ (.I(_4408_),
    .Z(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7751_ (.A1(_1416_),
    .A2(_2264_),
    .ZN(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7752_ (.A1(net50),
    .A2(_2941_),
    .B(_2308_),
    .C(_2942_),
    .ZN(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7753_ (.A1(_2940_),
    .A2(_2943_),
    .ZN(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7754_ (.A1(_1677_),
    .A2(_2937_),
    .B(_2938_),
    .C(_2944_),
    .ZN(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7755_ (.A1(net50),
    .A2(_2933_),
    .ZN(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7756_ (.A1(_2933_),
    .A2(_2945_),
    .B(_2946_),
    .C(_2437_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7757_ (.A1(_1616_),
    .A2(_2420_),
    .ZN(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7758_ (.A1(_2292_),
    .A2(_2418_),
    .B1(_2947_),
    .B2(_0940_),
    .ZN(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7759_ (.I(_2948_),
    .ZN(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7760_ (.A1(_2281_),
    .A2(_2148_),
    .ZN(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7761_ (.A1(_2145_),
    .A2(_1385_),
    .B(_2140_),
    .ZN(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7762_ (.A1(_2146_),
    .A2(_2950_),
    .A3(_2951_),
    .ZN(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7763_ (.A1(_4237_),
    .A2(_2145_),
    .A3(_2144_),
    .ZN(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7764_ (.A1(_2952_),
    .A2(_2953_),
    .ZN(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7765_ (.A1(_1631_),
    .A2(_2949_),
    .B(_2954_),
    .ZN(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7766_ (.I(_2272_),
    .Z(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7767_ (.I(_2956_),
    .Z(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7768_ (.A1(_1466_),
    .A2(_2957_),
    .B(_1183_),
    .ZN(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7769_ (.A1(_1447_),
    .A2(_2287_),
    .ZN(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7770_ (.I(_0924_),
    .Z(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7771_ (.I(_2314_),
    .Z(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7772_ (.A1(_2960_),
    .A2(_2961_),
    .B(_1378_),
    .ZN(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7773_ (.A1(_2238_),
    .A2(_2958_),
    .A3(_2959_),
    .A4(_2962_),
    .ZN(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _7774_ (.A1(_2258_),
    .A2(_2263_),
    .A3(_2955_),
    .A4(_2963_),
    .ZN(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7775_ (.I(_2964_),
    .ZN(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7776_ (.A1(_2303_),
    .A2(_2965_),
    .ZN(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7777_ (.I(_1456_),
    .Z(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7778_ (.A1(_2333_),
    .A2(_0929_),
    .ZN(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7779_ (.A1(net49),
    .A2(_2967_),
    .A3(_2968_),
    .ZN(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7780_ (.I(_2327_),
    .Z(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7781_ (.I(_2327_),
    .Z(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7782_ (.A1(_0948_),
    .A2(_2968_),
    .ZN(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7783_ (.A1(_2413_),
    .A2(_2972_),
    .ZN(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7784_ (.A1(net49),
    .A2(_2967_),
    .A3(_2971_),
    .A4(_2973_),
    .ZN(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7785_ (.A1(_2793_),
    .A2(_2970_),
    .B(_2974_),
    .ZN(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7786_ (.A1(net49),
    .A2(_2967_),
    .A3(_1436_),
    .ZN(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7787_ (.A1(_1633_),
    .A2(_2976_),
    .ZN(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7788_ (.A1(_2348_),
    .A2(_2975_),
    .B1(_2977_),
    .B2(_2223_),
    .ZN(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7789_ (.A1(_1488_),
    .A2(_2969_),
    .B1(_2978_),
    .B2(_1573_),
    .C(_2225_),
    .ZN(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7790_ (.A1(_2724_),
    .A2(_2979_),
    .ZN(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7791_ (.A1(net49),
    .A2(_2966_),
    .ZN(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7792_ (.I(_2436_),
    .Z(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7793_ (.A1(_2966_),
    .A2(_2980_),
    .B(_2981_),
    .C(_2982_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7794_ (.I(_2629_),
    .Z(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7795_ (.A1(_2983_),
    .A2(_1633_),
    .A3(_2132_),
    .ZN(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7796_ (.A1(_2587_),
    .A2(_2984_),
    .ZN(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _7797_ (.A1(_2233_),
    .A2(_2985_),
    .B(_2285_),
    .C(_2220_),
    .ZN(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7798_ (.A1(_2180_),
    .A2(_2309_),
    .ZN(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7799_ (.A1(_4452_),
    .A2(_2986_),
    .ZN(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7800_ (.A1(_2986_),
    .A2(_2987_),
    .B(_2988_),
    .C(_2982_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7801_ (.A1(_2182_),
    .A2(_2309_),
    .ZN(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7802_ (.A1(_4451_),
    .A2(_2986_),
    .ZN(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7803_ (.A1(_2986_),
    .A2(_2989_),
    .B(_2990_),
    .C(_2982_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7804_ (.I(_1351_),
    .Z(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7805_ (.A1(_2259_),
    .A2(_2261_),
    .ZN(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7806_ (.I(_0926_),
    .Z(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7807_ (.A1(_1659_),
    .A2(_4271_),
    .ZN(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7808_ (.A1(_1352_),
    .A2(_1565_),
    .B1(_2992_),
    .B2(_2993_),
    .C(_2994_),
    .ZN(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7809_ (.A1(_2991_),
    .A2(_4228_),
    .A3(_2992_),
    .B(_2995_),
    .ZN(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7810_ (.I(_2996_),
    .Z(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7811_ (.I(_2996_),
    .Z(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7812_ (.I(_1388_),
    .Z(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7813_ (.A1(_4353_),
    .A2(_2999_),
    .ZN(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7814_ (.A1(_2120_),
    .A2(_1638_),
    .B(_3000_),
    .ZN(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7815_ (.A1(_2998_),
    .A2(_3001_),
    .ZN(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7816_ (.A1(_4322_),
    .A2(_2997_),
    .B(_3002_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7817_ (.I(_1065_),
    .ZN(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7818_ (.I(_1395_),
    .Z(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7819_ (.A1(_1680_),
    .A2(_1639_),
    .ZN(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7820_ (.A1(_3003_),
    .A2(_3004_),
    .B(_3005_),
    .ZN(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7821_ (.I(_2996_),
    .Z(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7822_ (.I0(_3006_),
    .I1(\as2650.holding_reg[1] ),
    .S(_3007_),
    .Z(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7823_ (.I(_3008_),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7824_ (.I(_1577_),
    .Z(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7825_ (.I(_1394_),
    .Z(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7826_ (.A1(_0439_),
    .A2(_3010_),
    .ZN(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7827_ (.A1(_2167_),
    .A2(_3009_),
    .B(_3011_),
    .ZN(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7828_ (.I0(_3012_),
    .I1(\as2650.holding_reg[2] ),
    .S(_3007_),
    .Z(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7829_ (.I(_3013_),
    .Z(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7830_ (.I(_0543_),
    .ZN(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7831_ (.A1(_2171_),
    .A2(_2226_),
    .ZN(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7832_ (.A1(_3014_),
    .A2(_3004_),
    .B(_3015_),
    .ZN(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7833_ (.A1(_2998_),
    .A2(_3016_),
    .ZN(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7834_ (.A1(_0515_),
    .A2(_2997_),
    .B(_3017_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7835_ (.A1(_2176_),
    .A2(_2226_),
    .ZN(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7836_ (.A1(_1090_),
    .A2(_3009_),
    .B(_3018_),
    .ZN(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7837_ (.A1(_2998_),
    .A2(_3019_),
    .ZN(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7838_ (.A1(_0607_),
    .A2(_2997_),
    .B(_3020_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7839_ (.A1(_0783_),
    .A2(_2999_),
    .ZN(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7840_ (.A1(_2179_),
    .A2(_1624_),
    .B(_3021_),
    .ZN(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7841_ (.I0(_3022_),
    .I1(\as2650.holding_reg[5] ),
    .S(_3007_),
    .Z(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7842_ (.I(_3023_),
    .Z(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7843_ (.A1(_1689_),
    .A2(_1417_),
    .ZN(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7844_ (.A1(_1102_),
    .A2(_1634_),
    .ZN(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7845_ (.A1(\as2650.holding_reg[6] ),
    .A2(_2998_),
    .ZN(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7846_ (.A1(_2997_),
    .A2(_3024_),
    .A3(_3025_),
    .B(_3026_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7847_ (.A1(_2186_),
    .A2(_1417_),
    .B(_1625_),
    .ZN(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7848_ (.I0(_3027_),
    .I1(\as2650.holding_reg[7] ),
    .S(_3007_),
    .Z(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7849_ (.I(_3028_),
    .Z(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7850_ (.A1(_1634_),
    .A2(_2259_),
    .B(_2288_),
    .ZN(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7851_ (.A1(_2231_),
    .A2(_3029_),
    .Z(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7852_ (.I(_3030_),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7853_ (.A1(_2220_),
    .A2(_2230_),
    .ZN(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7854_ (.I(_3031_),
    .Z(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7855_ (.I(_2230_),
    .Z(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7856_ (.I(_2327_),
    .Z(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7857_ (.I(_2141_),
    .Z(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7858_ (.I(_3035_),
    .Z(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7859_ (.A1(_1154_),
    .A2(_2298_),
    .ZN(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7860_ (.I(_3037_),
    .Z(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7861_ (.I(_1442_),
    .Z(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7862_ (.A1(_3039_),
    .A2(_1659_),
    .A3(_2476_),
    .ZN(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7863_ (.A1(_3039_),
    .A2(_4254_),
    .B(_3036_),
    .ZN(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7864_ (.A1(_3036_),
    .A2(_3038_),
    .A3(_3040_),
    .B1(_3041_),
    .B2(_2527_),
    .ZN(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7865_ (.I(_3039_),
    .Z(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7866_ (.A1(_0926_),
    .A2(_1422_),
    .A3(_1402_),
    .A4(_1399_),
    .ZN(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7867_ (.A1(_3043_),
    .A2(_2412_),
    .B(_3044_),
    .ZN(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7868_ (.A1(_2339_),
    .A2(_2190_),
    .B(_3045_),
    .ZN(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7869_ (.I(_2209_),
    .Z(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7870_ (.A1(_2839_),
    .A2(_3042_),
    .B1(_3046_),
    .B2(_3047_),
    .ZN(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7871_ (.A1(_2993_),
    .A2(_3034_),
    .B1(_2225_),
    .B2(_3048_),
    .ZN(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7872_ (.A1(_2215_),
    .A2(_3049_),
    .ZN(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7873_ (.A1(_4444_),
    .A2(_4408_),
    .B1(_2361_),
    .B2(_2187_),
    .ZN(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7874_ (.A1(_2324_),
    .A2(_2941_),
    .B(_2368_),
    .ZN(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7875_ (.A1(_2531_),
    .A2(_2339_),
    .ZN(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7876_ (.A1(_3043_),
    .A2(_4267_),
    .B(_2200_),
    .C(_3053_),
    .ZN(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7877_ (.A1(_3051_),
    .A2(_3052_),
    .A3(_3054_),
    .ZN(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7878_ (.A1(_1634_),
    .A2(_1522_),
    .B(_2260_),
    .C(_3055_),
    .ZN(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7879_ (.A1(_3033_),
    .A2(_1474_),
    .A3(_3050_),
    .A4(_3056_),
    .ZN(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7880_ (.A1(_2993_),
    .A2(_3032_),
    .B(_3057_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7881_ (.I(_2991_),
    .Z(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7882_ (.A1(_2282_),
    .A2(_2283_),
    .A3(_3051_),
    .Z(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7883_ (.A1(_2748_),
    .A2(_3059_),
    .B(_3052_),
    .C(_2942_),
    .ZN(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7884_ (.A1(_3058_),
    .A2(_1522_),
    .B(_3060_),
    .ZN(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7885_ (.I(_2221_),
    .Z(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7886_ (.I(_3062_),
    .Z(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7887_ (.I(_1661_),
    .Z(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7888_ (.I(_1658_),
    .Z(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7889_ (.I(_3065_),
    .Z(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7890_ (.A1(_3066_),
    .A2(_2284_),
    .ZN(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7891_ (.I(_3035_),
    .Z(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7892_ (.I(_3068_),
    .Z(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7893_ (.A1(_3069_),
    .A2(_2264_),
    .ZN(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7894_ (.A1(_2971_),
    .A2(_2951_),
    .B(_2284_),
    .ZN(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7895_ (.A1(_3064_),
    .A2(_3038_),
    .B1(_3067_),
    .B2(_3070_),
    .C(_3071_),
    .ZN(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7896_ (.A1(_1633_),
    .A2(_3044_),
    .ZN(_3073_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7897_ (.A1(_2223_),
    .A2(_3067_),
    .A3(_3073_),
    .ZN(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7898_ (.A1(_3063_),
    .A2(_3072_),
    .B(_3074_),
    .C(_2588_),
    .ZN(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7899_ (.A1(_1632_),
    .A2(_3061_),
    .B(_3075_),
    .ZN(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7900_ (.A1(_0404_),
    .A2(_3032_),
    .B1(_3076_),
    .B2(_1031_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7901_ (.I(_2193_),
    .Z(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7902_ (.I(_3077_),
    .Z(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7903_ (.I(_2339_),
    .Z(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7904_ (.A1(_0927_),
    .A2(_2283_),
    .Z(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7905_ (.A1(_2967_),
    .A2(_1398_),
    .B(_3080_),
    .ZN(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7906_ (.A1(_2190_),
    .A2(_2198_),
    .B(_3081_),
    .ZN(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7907_ (.A1(_3079_),
    .A2(_2190_),
    .B(_3082_),
    .ZN(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7908_ (.A1(_3078_),
    .A2(_3083_),
    .ZN(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7909_ (.I(_2137_),
    .Z(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7910_ (.I(_3080_),
    .Z(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7911_ (.A1(_3079_),
    .A2(_2935_),
    .A3(_3085_),
    .A4(_3086_),
    .ZN(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7912_ (.I(_3035_),
    .Z(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7913_ (.I(_3088_),
    .Z(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7914_ (.A1(_3043_),
    .A2(_2145_),
    .B(_3089_),
    .C(_3086_),
    .ZN(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7915_ (.I(_2344_),
    .Z(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7916_ (.I(_3091_),
    .Z(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7917_ (.A1(_0406_),
    .A2(_3092_),
    .B1(_2527_),
    .B2(_3089_),
    .C(_3047_),
    .ZN(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7918_ (.A1(_3087_),
    .A2(_3090_),
    .A3(_3093_),
    .ZN(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7919_ (.I(_2939_),
    .Z(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7920_ (.A1(_3084_),
    .A2(_3094_),
    .B(_3095_),
    .ZN(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7921_ (.I(_1420_),
    .Z(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _7922_ (.A1(_1349_),
    .A2(_3097_),
    .A3(_0334_),
    .A4(_1471_),
    .ZN(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7923_ (.A1(_0409_),
    .A2(_3086_),
    .B(_3098_),
    .C(_2280_),
    .ZN(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7924_ (.I(_2235_),
    .Z(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7925_ (.I(_3100_),
    .Z(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7926_ (.A1(_3101_),
    .A2(_2382_),
    .ZN(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7927_ (.A1(_3086_),
    .A2(_3102_),
    .B(_0963_),
    .ZN(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7928_ (.A1(_3096_),
    .A2(_3099_),
    .A3(_3103_),
    .B1(_3031_),
    .B2(_0927_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7929_ (.I(_2220_),
    .Z(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7930_ (.A1(_4238_),
    .A2(_4120_),
    .A3(_0943_),
    .A4(_3039_),
    .ZN(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7931_ (.A1(_0927_),
    .A2(_2283_),
    .B(_4188_),
    .ZN(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7932_ (.A1(_3105_),
    .A2(_3106_),
    .ZN(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7933_ (.A1(_4444_),
    .A2(_2941_),
    .A3(_2922_),
    .ZN(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7934_ (.A1(_2186_),
    .A2(_2941_),
    .A3(_2748_),
    .ZN(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7935_ (.A1(_3107_),
    .A2(_3108_),
    .A3(_3109_),
    .ZN(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7936_ (.A1(_1573_),
    .A2(_2264_),
    .A3(_2200_),
    .ZN(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7937_ (.A1(_3110_),
    .A2(_3111_),
    .ZN(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7938_ (.A1(_2332_),
    .A2(_0409_),
    .A3(_1660_),
    .B(_2947_),
    .ZN(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7939_ (.I(_2222_),
    .Z(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7940_ (.A1(_2217_),
    .A2(_1660_),
    .A3(_2968_),
    .B(_3085_),
    .ZN(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7941_ (.A1(_3114_),
    .A2(_3115_),
    .B(_3107_),
    .C(_2917_),
    .ZN(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7942_ (.A1(_2797_),
    .A2(_3113_),
    .B(_3116_),
    .C(_3104_),
    .ZN(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7943_ (.I(_1427_),
    .Z(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7944_ (.A1(_3104_),
    .A2(_4188_),
    .B1(_3112_),
    .B2(_3117_),
    .C(_3118_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7945_ (.I(\as2650.cycle[4] ),
    .Z(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7946_ (.A1(_2199_),
    .A2(_3105_),
    .ZN(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7947_ (.A1(_3119_),
    .A2(_3120_),
    .B(_2852_),
    .ZN(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7948_ (.A1(_3119_),
    .A2(_3120_),
    .B(_3121_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7949_ (.I(_1427_),
    .Z(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7950_ (.I(_3122_),
    .Z(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7951_ (.A1(_3119_),
    .A2(_3120_),
    .ZN(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7952_ (.A1(_4121_),
    .A2(_3124_),
    .Z(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7953_ (.A1(_3123_),
    .A2(_3125_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7954_ (.I(_2917_),
    .Z(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7955_ (.I(_4187_),
    .Z(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7956_ (.I(_3127_),
    .Z(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7957_ (.A1(_1682_),
    .A2(_3128_),
    .B(_2918_),
    .C(_2922_),
    .ZN(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7958_ (.A1(_4121_),
    .A2(_3119_),
    .ZN(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7959_ (.A1(_3105_),
    .A2(_3130_),
    .Z(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7960_ (.A1(_2562_),
    .A2(_3131_),
    .Z(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7961_ (.A1(_2562_),
    .A2(_3131_),
    .ZN(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7962_ (.A1(_3132_),
    .A2(_3133_),
    .ZN(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7963_ (.A1(_4444_),
    .A2(_3126_),
    .B(_3134_),
    .ZN(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7964_ (.A1(_3126_),
    .A2(_3129_),
    .B(_3135_),
    .C(_3104_),
    .ZN(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7965_ (.A1(_3104_),
    .A2(_2562_),
    .B(_3118_),
    .C(_3136_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7966_ (.A1(_1475_),
    .A2(_1350_),
    .ZN(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7967_ (.I(_3137_),
    .Z(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7968_ (.I(_2361_),
    .Z(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7969_ (.A1(_3004_),
    .A2(_3139_),
    .A3(_2748_),
    .B(_3126_),
    .ZN(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7970_ (.A1(_4443_),
    .A2(_3132_),
    .Z(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7971_ (.A1(_3138_),
    .A2(_3126_),
    .B1(_3140_),
    .B2(_3141_),
    .ZN(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7972_ (.A1(_4443_),
    .A2(_3032_),
    .B1(_3142_),
    .B2(_1031_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7973_ (.I(\as2650.psu[7] ),
    .ZN(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7974_ (.A1(_1691_),
    .A2(_1413_),
    .ZN(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7975_ (.A1(\as2650.psu[7] ),
    .A2(_1691_),
    .B(_3144_),
    .ZN(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7976_ (.A1(net4),
    .A2(_1404_),
    .ZN(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7977_ (.A1(_0861_),
    .A2(_1467_),
    .B(_3097_),
    .ZN(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7978_ (.A1(_1457_),
    .A2(_3145_),
    .B1(_3146_),
    .B2(_3147_),
    .ZN(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _7979_ (.A1(net4),
    .A2(_3004_),
    .A3(_1457_),
    .Z(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7980_ (.A1(_0963_),
    .A2(_3148_),
    .A3(_3149_),
    .ZN(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7981_ (.A1(_3143_),
    .A2(_3032_),
    .B(_3150_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7982_ (.A1(_4443_),
    .A2(_2122_),
    .B(_1455_),
    .C(_2968_),
    .ZN(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7983_ (.A1(_2143_),
    .A2(_2473_),
    .B(_2191_),
    .C(_0923_),
    .ZN(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7984_ (.A1(_1511_),
    .A2(_3152_),
    .ZN(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7985_ (.A1(_1523_),
    .A2(_3151_),
    .B(_3153_),
    .ZN(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7986_ (.A1(_2251_),
    .A2(_2271_),
    .A3(_2921_),
    .ZN(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7987_ (.A1(_1390_),
    .A2(_2256_),
    .B1(_2474_),
    .B2(_2141_),
    .C(_3155_),
    .ZN(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7988_ (.A1(_1350_),
    .A2(_1521_),
    .ZN(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7989_ (.A1(_1357_),
    .A2(_3157_),
    .B(_2287_),
    .ZN(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7990_ (.A1(_2267_),
    .A2(_3154_),
    .A3(_3156_),
    .A4(_3158_),
    .Z(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7991_ (.A1(_2255_),
    .A2(_2262_),
    .ZN(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7992_ (.A1(_2143_),
    .A2(_2950_),
    .A3(_2972_),
    .B(_2266_),
    .ZN(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7993_ (.A1(_4115_),
    .A2(_2302_),
    .A3(_2926_),
    .Z(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7994_ (.A1(_2280_),
    .A2(_2285_),
    .B(_2954_),
    .C(_3162_),
    .ZN(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7995_ (.A1(_3160_),
    .A2(_3161_),
    .A3(_3163_),
    .ZN(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7996_ (.A1(_3159_),
    .A2(_3164_),
    .ZN(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7997_ (.I(_3165_),
    .Z(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7998_ (.I(_3166_),
    .Z(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7999_ (.I(_2939_),
    .Z(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8000_ (.A1(_2161_),
    .A2(_0408_),
    .ZN(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8001_ (.A1(_2336_),
    .A2(_3169_),
    .B(_3065_),
    .ZN(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8002_ (.I(_0901_),
    .Z(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8003_ (.A1(_1057_),
    .A2(_3171_),
    .ZN(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8004_ (.A1(_1544_),
    .A2(_2325_),
    .B(_3172_),
    .ZN(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8005_ (.A1(_1057_),
    .A2(_0938_),
    .ZN(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8006_ (.A1(_1682_),
    .A2(_3173_),
    .B(_3174_),
    .C(_1456_),
    .ZN(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8007_ (.A1(_1055_),
    .A2(_4197_),
    .ZN(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8008_ (.A1(_3174_),
    .A2(_3176_),
    .ZN(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8009_ (.I0(_3177_),
    .I1(_2310_),
    .S(_2297_),
    .Z(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8010_ (.A1(_2296_),
    .A2(_3177_),
    .ZN(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8011_ (.A1(_1057_),
    .A2(_2296_),
    .B(_3179_),
    .C(_4183_),
    .ZN(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8012_ (.A1(_4183_),
    .A2(_3178_),
    .B(_3180_),
    .C(_1351_),
    .ZN(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8013_ (.I(_0948_),
    .Z(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8014_ (.I(_3182_),
    .Z(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _8015_ (.A1(_3170_),
    .A2(_3175_),
    .A3(_3181_),
    .B(_3183_),
    .ZN(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8016_ (.A1(_2340_),
    .A2(_4302_),
    .ZN(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8017_ (.A1(_1203_),
    .A2(_3185_),
    .Z(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8018_ (.A1(_2311_),
    .A2(_1659_),
    .ZN(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8019_ (.A1(_2412_),
    .A2(_3186_),
    .B(_3187_),
    .C(_3036_),
    .ZN(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8020_ (.A1(_2970_),
    .A2(_3184_),
    .A3(_3188_),
    .ZN(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8021_ (.I(_0940_),
    .Z(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8022_ (.I(_3190_),
    .Z(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8023_ (.A1(_2311_),
    .A2(_3127_),
    .B1(_2873_),
    .B2(_3173_),
    .C(_3191_),
    .ZN(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8024_ (.A1(_3189_),
    .A2(_3192_),
    .ZN(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8025_ (.A1(_4471_),
    .A2(_4483_),
    .ZN(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8026_ (.I(_3194_),
    .Z(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8027_ (.I(_3195_),
    .Z(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8028_ (.A1(_0383_),
    .A2(\as2650.stack[1][0] ),
    .B1(\as2650.stack[0][0] ),
    .B2(_0386_),
    .ZN(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8029_ (.A1(_3196_),
    .A2(_3197_),
    .Z(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8030_ (.I(_0376_),
    .Z(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8031_ (.I(_3199_),
    .Z(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8032_ (.A1(_0918_),
    .A2(\as2650.stack[3][0] ),
    .B1(\as2650.stack[2][0] ),
    .B2(_3200_),
    .C(_4488_),
    .ZN(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8033_ (.I(_0380_),
    .Z(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8034_ (.I(\as2650.stack[6][0] ),
    .ZN(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8035_ (.I(_3194_),
    .Z(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8036_ (.I(_0379_),
    .Z(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8037_ (.A1(_0493_),
    .A2(\as2650.stack[5][0] ),
    .B1(\as2650.stack[4][0] ),
    .B2(_3205_),
    .ZN(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8038_ (.A1(_3203_),
    .A2(_4472_),
    .B1(_3204_),
    .B2(_3206_),
    .ZN(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8039_ (.A1(\as2650.stack[7][0] ),
    .A2(_3202_),
    .B(_0501_),
    .C(_3207_),
    .ZN(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8040_ (.A1(_3198_),
    .A2(_3201_),
    .B(_3208_),
    .ZN(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8041_ (.I(_3100_),
    .Z(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8042_ (.A1(_1058_),
    .A2(_3077_),
    .B1(_3209_),
    .B2(_3210_),
    .ZN(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8043_ (.I(_2244_),
    .Z(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8044_ (.A1(_3193_),
    .A2(_3211_),
    .B(_3212_),
    .ZN(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8045_ (.I(_3165_),
    .Z(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8046_ (.A1(_1058_),
    .A2(_3168_),
    .B(_3213_),
    .C(_3214_),
    .ZN(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8047_ (.A1(_1058_),
    .A2(_3167_),
    .B(_3215_),
    .C(_2982_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8048_ (.A1(_2380_),
    .A2(_1056_),
    .Z(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8049_ (.I(_3216_),
    .Z(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8050_ (.I(_2193_),
    .Z(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8051_ (.A1(_3218_),
    .A2(_3217_),
    .ZN(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8052_ (.A1(net6),
    .A2(_4302_),
    .ZN(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8053_ (.A1(_0351_),
    .A2(_4380_),
    .A3(_3220_),
    .Z(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8054_ (.A1(_0352_),
    .A2(_2338_),
    .B(_2216_),
    .ZN(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8055_ (.A1(_2596_),
    .A2(_3221_),
    .B(_3222_),
    .ZN(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8056_ (.I(_2420_),
    .Z(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8057_ (.A1(_2184_),
    .A2(_2425_),
    .ZN(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8058_ (.A1(_2380_),
    .A2(_2604_),
    .B(_3225_),
    .ZN(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8059_ (.A1(_2803_),
    .A2(_2130_),
    .B(_2141_),
    .ZN(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8060_ (.A1(_0352_),
    .A2(_2338_),
    .B1(_2417_),
    .B2(_3216_),
    .C(_3227_),
    .ZN(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8061_ (.A1(_3224_),
    .A2(_3226_),
    .B(_3228_),
    .ZN(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8062_ (.A1(_3036_),
    .A2(_3223_),
    .B(_3229_),
    .C(_1577_),
    .ZN(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8063_ (.I(_2299_),
    .Z(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8064_ (.A1(_1068_),
    .A2(_3176_),
    .Z(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _8065_ (.A1(_3035_),
    .A2(_3037_),
    .B(_3065_),
    .ZN(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _8066_ (.A1(_3068_),
    .A2(_3231_),
    .A3(_3232_),
    .B1(_3233_),
    .B2(_3217_),
    .ZN(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8067_ (.A1(_3230_),
    .A2(_3234_),
    .B(_2971_),
    .ZN(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8068_ (.A1(_3137_),
    .A2(_3217_),
    .ZN(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8069_ (.A1(_2313_),
    .A2(_3226_),
    .B(_3236_),
    .C(_3190_),
    .ZN(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8070_ (.I(_0379_),
    .Z(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8071_ (.A1(_0493_),
    .A2(\as2650.stack[1][1] ),
    .B1(\as2650.stack[0][1] ),
    .B2(_3238_),
    .ZN(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8072_ (.A1(_3204_),
    .A2(_3239_),
    .Z(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8073_ (.I(_4487_),
    .Z(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8074_ (.A1(_1590_),
    .A2(\as2650.stack[3][1] ),
    .B1(\as2650.stack[2][1] ),
    .B2(_0377_),
    .C(_3241_),
    .ZN(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8075_ (.I(_0380_),
    .Z(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8076_ (.I(\as2650.stack[6][1] ),
    .ZN(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8077_ (.I(_4469_),
    .Z(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8078_ (.A1(_3245_),
    .A2(\as2650.stack[5][1] ),
    .B1(\as2650.stack[4][1] ),
    .B2(_0385_),
    .ZN(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8079_ (.A1(_3244_),
    .A2(_4471_),
    .B1(_3195_),
    .B2(_3246_),
    .ZN(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8080_ (.A1(\as2650.stack[7][1] ),
    .A2(_3243_),
    .B(_4497_),
    .C(_3247_),
    .ZN(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8081_ (.A1(_3240_),
    .A2(_3242_),
    .B(_3248_),
    .ZN(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8082_ (.A1(_3235_),
    .A2(_3237_),
    .B1(_3249_),
    .B2(_3210_),
    .ZN(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8083_ (.I(_2244_),
    .Z(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8084_ (.A1(_3219_),
    .A2(_3250_),
    .B(_3251_),
    .ZN(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8085_ (.A1(_3168_),
    .A2(_3217_),
    .B(_3252_),
    .C(_3214_),
    .ZN(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8086_ (.I(_2436_),
    .Z(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8087_ (.A1(_1068_),
    .A2(_3167_),
    .B(_3253_),
    .C(_3254_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8088_ (.I(_2245_),
    .Z(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8089_ (.A1(_1066_),
    .A2(_1056_),
    .ZN(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8090_ (.A1(_1074_),
    .A2(_3256_),
    .ZN(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8091_ (.A1(_1074_),
    .A2(_3256_),
    .Z(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8092_ (.A1(_1074_),
    .A2(_1616_),
    .ZN(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8093_ (.A1(_1544_),
    .A2(_2482_),
    .B(_3259_),
    .ZN(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8094_ (.A1(_2531_),
    .A2(_3260_),
    .ZN(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8095_ (.A1(_2615_),
    .A2(_3258_),
    .B(_3261_),
    .C(_3091_),
    .ZN(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8096_ (.I(_2299_),
    .Z(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8097_ (.A1(_1067_),
    .A2(_3176_),
    .ZN(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8098_ (.A1(_1075_),
    .A2(_3264_),
    .Z(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8099_ (.I(_3037_),
    .Z(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8100_ (.A1(_3224_),
    .A2(_3260_),
    .ZN(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8101_ (.A1(_2168_),
    .A2(_2197_),
    .ZN(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8102_ (.A1(_1155_),
    .A2(_3268_),
    .ZN(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _8103_ (.A1(_1552_),
    .A2(_2778_),
    .B1(_2961_),
    .B2(_3257_),
    .C(_3269_),
    .ZN(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8104_ (.A1(_3266_),
    .A2(_3258_),
    .B1(_3267_),
    .B2(_3270_),
    .C(_3068_),
    .ZN(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8105_ (.A1(_3263_),
    .A2(_3265_),
    .B(_3271_),
    .ZN(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8106_ (.I(_1443_),
    .Z(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8107_ (.I(_3273_),
    .Z(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8108_ (.A1(_0453_),
    .A2(_0340_),
    .Z(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8109_ (.A1(_0349_),
    .A2(_4380_),
    .ZN(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8110_ (.A1(_2440_),
    .A2(_4380_),
    .ZN(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8111_ (.A1(_3220_),
    .A2(_3276_),
    .B(_3277_),
    .ZN(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8112_ (.A1(_3275_),
    .A2(_3278_),
    .ZN(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8113_ (.I(_0407_),
    .Z(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8114_ (.A1(_1552_),
    .A2(_3280_),
    .ZN(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8115_ (.A1(_2596_),
    .A2(_3279_),
    .B(_3281_),
    .C(_3273_),
    .ZN(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8116_ (.A1(_3274_),
    .A2(_3257_),
    .B(_3282_),
    .C(_3069_),
    .ZN(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8117_ (.A1(_3034_),
    .A2(_3272_),
    .A3(_3283_),
    .ZN(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8118_ (.A1(_3262_),
    .A2(_3284_),
    .ZN(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8119_ (.A1(_3063_),
    .A2(_3285_),
    .ZN(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8120_ (.I(_3077_),
    .Z(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8121_ (.I(\as2650.stack[6][2] ),
    .ZN(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8122_ (.A1(_0493_),
    .A2(\as2650.stack[5][2] ),
    .B1(\as2650.stack[4][2] ),
    .B2(_3205_),
    .ZN(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8123_ (.A1(_3288_),
    .A2(_4472_),
    .B1(_3204_),
    .B2(_3289_),
    .ZN(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8124_ (.A1(\as2650.stack[7][2] ),
    .A2(_3243_),
    .B(_0501_),
    .C(_3290_),
    .ZN(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8125_ (.I(\as2650.stack[2][2] ),
    .ZN(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8126_ (.A1(_3245_),
    .A2(\as2650.stack[1][2] ),
    .B1(\as2650.stack[0][2] ),
    .B2(_3205_),
    .ZN(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8127_ (.A1(_3292_),
    .A2(_4472_),
    .B1(_3204_),
    .B2(_3293_),
    .ZN(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8128_ (.A1(\as2650.stack[3][2] ),
    .A2(_3243_),
    .B(_3241_),
    .C(_3294_),
    .ZN(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8129_ (.A1(_3291_),
    .A2(_3295_),
    .ZN(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8130_ (.I(_3296_),
    .ZN(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8131_ (.A1(_3287_),
    .A2(_3258_),
    .B1(_3297_),
    .B2(_3101_),
    .C(_2940_),
    .ZN(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8132_ (.I(_3165_),
    .Z(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8133_ (.I(_3299_),
    .Z(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8134_ (.A1(_3255_),
    .A2(_3257_),
    .B1(_3286_),
    .B2(_3298_),
    .C(_3300_),
    .ZN(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8135_ (.A1(_3159_),
    .A2(_3164_),
    .Z(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8136_ (.I(_3302_),
    .Z(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8137_ (.A1(_1076_),
    .A2(_3303_),
    .B(_3033_),
    .ZN(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8138_ (.A1(_3301_),
    .A2(_3304_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _8139_ (.A1(\as2650.pc[2] ),
    .A2(\as2650.pc[1] ),
    .A3(\as2650.pc[0] ),
    .ZN(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8140_ (.A1(_1083_),
    .A2(_3305_),
    .Z(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8141_ (.A1(_3218_),
    .A2(_3306_),
    .ZN(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _8142_ (.A1(_2491_),
    .A2(_1073_),
    .A3(_3264_),
    .Z(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8143_ (.A1(_1075_),
    .A2(_3264_),
    .B(_2492_),
    .ZN(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8144_ (.A1(_1465_),
    .A2(_2298_),
    .Z(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8145_ (.A1(_3308_),
    .A2(_3309_),
    .B(_3310_),
    .ZN(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8146_ (.A1(_2492_),
    .A2(_3305_),
    .Z(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8147_ (.A1(_3266_),
    .A2(_3312_),
    .ZN(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8148_ (.A1(_1083_),
    .A2(_0902_),
    .ZN(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8149_ (.A1(_3171_),
    .A2(_2522_),
    .B(_3314_),
    .ZN(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _8150_ (.A1(_1555_),
    .A2(_2340_),
    .B1(_2197_),
    .B2(_2172_),
    .C(_1465_),
    .ZN(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8151_ (.A1(_2418_),
    .A2(_3312_),
    .B1(_3315_),
    .B2(_3085_),
    .C(_3316_),
    .ZN(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8152_ (.A1(_2934_),
    .A2(_3311_),
    .A3(_3313_),
    .A4(_3317_),
    .ZN(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8153_ (.A1(_0453_),
    .A2(_0340_),
    .Z(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8154_ (.A1(_3275_),
    .A2(_3278_),
    .B(_3319_),
    .ZN(_3320_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8155_ (.A1(_1554_),
    .A2(_0446_),
    .A3(_3320_),
    .Z(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8156_ (.A1(_1555_),
    .A2(_3280_),
    .ZN(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8157_ (.A1(_2596_),
    .A2(_3321_),
    .B(_3322_),
    .C(_1443_),
    .ZN(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8158_ (.A1(_2841_),
    .A2(_3306_),
    .B(_3323_),
    .C(_3088_),
    .ZN(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8159_ (.A1(_2971_),
    .A2(_3318_),
    .A3(_3324_),
    .ZN(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8160_ (.A1(_3127_),
    .A2(_3312_),
    .B1(_3315_),
    .B2(_2313_),
    .C(_3190_),
    .ZN(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8161_ (.I(_3195_),
    .Z(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8162_ (.I(_0385_),
    .Z(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8163_ (.A1(_0494_),
    .A2(\as2650.stack[1][3] ),
    .B1(\as2650.stack[0][3] ),
    .B2(_3328_),
    .ZN(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8164_ (.A1(_3327_),
    .A2(_3329_),
    .Z(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8165_ (.I(_0377_),
    .Z(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8166_ (.A1(_0919_),
    .A2(\as2650.stack[3][3] ),
    .B1(\as2650.stack[2][3] ),
    .B2(_3331_),
    .C(_4488_),
    .ZN(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8167_ (.I(\as2650.stack[6][3] ),
    .ZN(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8168_ (.A1(_0383_),
    .A2(\as2650.stack[5][3] ),
    .B1(\as2650.stack[4][3] ),
    .B2(_3328_),
    .ZN(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8169_ (.A1(_3333_),
    .A2(_4475_),
    .B1(_3327_),
    .B2(_3334_),
    .ZN(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8170_ (.A1(\as2650.stack[7][3] ),
    .A2(_3202_),
    .B(_4498_),
    .C(_3335_),
    .ZN(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8171_ (.A1(_3330_),
    .A2(_3332_),
    .B(_3336_),
    .ZN(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8172_ (.A1(_3325_),
    .A2(_3326_),
    .B1(_3337_),
    .B2(_3210_),
    .ZN(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8173_ (.A1(_3307_),
    .A2(_3338_),
    .B(_3251_),
    .ZN(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8174_ (.A1(_3168_),
    .A2(_3306_),
    .B(_3339_),
    .C(_3214_),
    .ZN(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8175_ (.A1(_1084_),
    .A2(_3167_),
    .B(_3340_),
    .C(_3254_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8176_ (.I(_3214_),
    .Z(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8177_ (.A1(_2587_),
    .A2(_2381_),
    .ZN(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8178_ (.I(_3342_),
    .Z(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8179_ (.A1(_1083_),
    .A2(_3305_),
    .ZN(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8180_ (.A1(_2540_),
    .A2(_3344_),
    .Z(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8181_ (.I(_3345_),
    .Z(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8182_ (.I(_3233_),
    .Z(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8183_ (.A1(_2541_),
    .A2(_3308_),
    .Z(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8184_ (.A1(_1288_),
    .A2(_0407_),
    .Z(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8185_ (.A1(_2144_),
    .A2(_3349_),
    .ZN(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8186_ (.A1(_0676_),
    .A2(_0547_),
    .Z(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8187_ (.A1(_0554_),
    .A2(_0446_),
    .ZN(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8188_ (.A1(_0554_),
    .A2(_0446_),
    .ZN(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8189_ (.A1(_3352_),
    .A2(_3320_),
    .B(_3353_),
    .ZN(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8190_ (.A1(_3351_),
    .A2(_3354_),
    .B(_4256_),
    .ZN(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8191_ (.A1(_3351_),
    .A2(_3354_),
    .B(_3355_),
    .ZN(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8192_ (.I(_2314_),
    .Z(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8193_ (.A1(_2541_),
    .A2(_1543_),
    .ZN(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8194_ (.A1(_0902_),
    .A2(_2582_),
    .B(_3358_),
    .ZN(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8195_ (.I(_0932_),
    .Z(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8196_ (.A1(_0677_),
    .A2(_2206_),
    .B1(_2130_),
    .B2(\as2650.addr_buff[4] ),
    .ZN(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8197_ (.A1(_2150_),
    .A2(_3361_),
    .ZN(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _8198_ (.A1(_3357_),
    .A2(_3345_),
    .B1(_3359_),
    .B2(_3360_),
    .C(_3362_),
    .ZN(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8199_ (.A1(_3350_),
    .A2(_3356_),
    .B(_3363_),
    .ZN(_3364_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _8200_ (.A1(_3088_),
    .A2(_3231_),
    .A3(_3348_),
    .B1(_3364_),
    .B2(_1416_),
    .ZN(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8201_ (.A1(_3137_),
    .A2(_3346_),
    .B1(_3359_),
    .B2(_2572_),
    .C(_2837_),
    .ZN(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8202_ (.A1(_2970_),
    .A2(_3365_),
    .B(_3366_),
    .ZN(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8203_ (.A1(_3347_),
    .A2(_3346_),
    .B1(_3367_),
    .B2(_2245_),
    .ZN(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8204_ (.I(_3100_),
    .Z(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8205_ (.A1(_1582_),
    .A2(\as2650.stack[5][4] ),
    .B1(\as2650.stack[4][4] ),
    .B2(_3238_),
    .ZN(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8206_ (.A1(_3196_),
    .A2(_3370_),
    .Z(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _8207_ (.A1(\as2650.stack[6][4] ),
    .A2(_3200_),
    .B1(_3243_),
    .B2(\as2650.stack[7][4] ),
    .C(_4497_),
    .ZN(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8208_ (.A1(_1582_),
    .A2(\as2650.stack[1][4] ),
    .B1(\as2650.stack[0][4] ),
    .B2(_3238_),
    .ZN(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8209_ (.A1(_3196_),
    .A2(_3373_),
    .Z(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _8210_ (.A1(_1590_),
    .A2(\as2650.stack[3][4] ),
    .B1(\as2650.stack[2][4] ),
    .B2(_0377_),
    .C(_3241_),
    .ZN(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _8211_ (.A1(_3371_),
    .A2(_3372_),
    .B1(_3374_),
    .B2(_3375_),
    .ZN(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8212_ (.A1(_3369_),
    .A2(_3376_),
    .ZN(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8213_ (.A1(_3368_),
    .A2(_3377_),
    .ZN(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8214_ (.A1(_3343_),
    .A2(_3346_),
    .B(_3378_),
    .ZN(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8215_ (.A1(_3078_),
    .A2(_3346_),
    .B(_3166_),
    .ZN(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8216_ (.A1(_1091_),
    .A2(_3341_),
    .B1(_3379_),
    .B2(_3380_),
    .C(_3122_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8217_ (.A1(_1091_),
    .A2(_1082_),
    .A3(_3305_),
    .ZN(_3381_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8218_ (.A1(_2594_),
    .A2(_3381_),
    .Z(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8219_ (.A1(_1097_),
    .A2(_3381_),
    .Z(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8220_ (.A1(_3065_),
    .A2(_3182_),
    .ZN(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8221_ (.A1(_0674_),
    .A2(_0547_),
    .Z(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8222_ (.A1(_0674_),
    .A2(_0547_),
    .Z(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8223_ (.A1(_3385_),
    .A2(_3354_),
    .B(_3386_),
    .ZN(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8224_ (.A1(_0758_),
    .A2(_0652_),
    .A3(_3387_),
    .Z(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8225_ (.A1(_1410_),
    .A2(_2475_),
    .ZN(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8226_ (.A1(_2476_),
    .A2(_3388_),
    .B(_3389_),
    .ZN(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8227_ (.A1(_2540_),
    .A2(_3308_),
    .ZN(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8228_ (.A1(_2595_),
    .A2(_3391_),
    .Z(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8229_ (.A1(_1581_),
    .A2(_2611_),
    .ZN(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8230_ (.A1(_2595_),
    .A2(_2184_),
    .B(_3393_),
    .ZN(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8231_ (.A1(_3360_),
    .A2(_3394_),
    .Z(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8232_ (.A1(_2180_),
    .A2(_0407_),
    .ZN(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8233_ (.A1(_1585_),
    .A2(_3280_),
    .B(_3396_),
    .C(_1373_),
    .ZN(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8234_ (.A1(_2418_),
    .A2(_3382_),
    .B(_3397_),
    .C(_1419_),
    .ZN(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8235_ (.A1(_2299_),
    .A2(_3392_),
    .B1(_3395_),
    .B2(_3398_),
    .ZN(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8236_ (.A1(_3384_),
    .A2(_3390_),
    .B1(_3399_),
    .B2(_2934_),
    .C(_3091_),
    .ZN(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8237_ (.A1(_3233_),
    .A2(_3383_),
    .B(_3400_),
    .ZN(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8238_ (.A1(_3127_),
    .A2(_3383_),
    .B1(_3394_),
    .B2(_2873_),
    .C(_3190_),
    .ZN(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8239_ (.A1(_3401_),
    .A2(_3402_),
    .ZN(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8240_ (.A1(_3205_),
    .A2(\as2650.stack[1][5] ),
    .B1(\as2650.stack[0][5] ),
    .B2(_3245_),
    .ZN(_3404_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8241_ (.A1(_3199_),
    .A2(_3404_),
    .Z(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8242_ (.A1(_1590_),
    .A2(\as2650.stack[3][5] ),
    .B1(\as2650.stack[2][5] ),
    .B2(_3199_),
    .C(_4487_),
    .ZN(_3406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8243_ (.A1(_3245_),
    .A2(\as2650.stack[5][5] ),
    .B1(\as2650.stack[4][5] ),
    .B2(_0385_),
    .ZN(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8244_ (.A1(_3195_),
    .A2(_3407_),
    .Z(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8245_ (.A1(\as2650.stack[6][5] ),
    .A2(_3199_),
    .B1(_0380_),
    .B2(\as2650.stack[7][5] ),
    .C(_4497_),
    .ZN(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8246_ (.A1(_3405_),
    .A2(_3406_),
    .B1(_3408_),
    .B2(_3409_),
    .ZN(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8247_ (.A1(_3218_),
    .A2(_3382_),
    .B1(_3410_),
    .B2(_3210_),
    .ZN(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8248_ (.A1(_3403_),
    .A2(_3411_),
    .B(_3251_),
    .ZN(_3412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8249_ (.A1(_3168_),
    .A2(_3382_),
    .B(_3412_),
    .C(_3299_),
    .ZN(_3413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8250_ (.A1(_1097_),
    .A2(_3167_),
    .B(_3413_),
    .C(_3254_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8251_ (.A1(_2594_),
    .A2(_3381_),
    .ZN(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8252_ (.A1(_1105_),
    .A2(_3414_),
    .Z(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8253_ (.I(_3415_),
    .Z(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8254_ (.A1(_1103_),
    .A2(_3171_),
    .ZN(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8255_ (.A1(_1621_),
    .A2(_2681_),
    .B(_3417_),
    .ZN(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8256_ (.I(_3360_),
    .Z(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8257_ (.A1(_1525_),
    .A2(_2236_),
    .ZN(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8258_ (.A1(_2182_),
    .A2(_3280_),
    .ZN(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8259_ (.A1(_3420_),
    .A2(_3421_),
    .B(_2601_),
    .ZN(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8260_ (.A1(_2961_),
    .A2(_3415_),
    .B1(_3418_),
    .B2(_3419_),
    .C(_3422_),
    .ZN(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8261_ (.A1(_2594_),
    .A2(_2539_),
    .A3(_3308_),
    .ZN(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8262_ (.A1(_2647_),
    .A2(_3424_),
    .Z(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8263_ (.A1(_3010_),
    .A2(_3423_),
    .B1(_3425_),
    .B2(_3231_),
    .C(_3183_),
    .ZN(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8264_ (.A1(_3038_),
    .A2(_3416_),
    .B(_3426_),
    .ZN(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8265_ (.A1(_2606_),
    .A2(_0652_),
    .ZN(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8266_ (.A1(_2606_),
    .A2(_0652_),
    .ZN(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8267_ (.A1(_3428_),
    .A2(_3387_),
    .B(_3429_),
    .ZN(_3430_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _8268_ (.A1(_0833_),
    .A2(_0747_),
    .A3(_3430_),
    .ZN(_3431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8269_ (.A1(_1559_),
    .A2(_2528_),
    .B(_3273_),
    .ZN(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8270_ (.A1(_2677_),
    .A2(_3431_),
    .B(_3432_),
    .ZN(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8271_ (.A1(_3066_),
    .A2(_3415_),
    .B(_3433_),
    .C(_2935_),
    .ZN(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8272_ (.A1(_3128_),
    .A2(_3416_),
    .B1(_3418_),
    .B2(_2873_),
    .C(_3191_),
    .ZN(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _8273_ (.A1(_3092_),
    .A2(_3427_),
    .A3(_3434_),
    .B(_3435_),
    .ZN(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8274_ (.A1(\as2650.stack[6][6] ),
    .A2(_3331_),
    .B1(_3202_),
    .B2(\as2650.stack[7][6] ),
    .ZN(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8275_ (.I0(\as2650.stack[5][6] ),
    .I1(\as2650.stack[4][6] ),
    .S(_4468_),
    .Z(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8276_ (.A1(_0381_),
    .A2(_3438_),
    .B(_4498_),
    .ZN(_3439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8277_ (.A1(_0494_),
    .A2(\as2650.stack[1][6] ),
    .B1(\as2650.stack[0][6] ),
    .B2(_3328_),
    .ZN(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8278_ (.A1(_3327_),
    .A2(_3440_),
    .Z(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8279_ (.A1(_0918_),
    .A2(\as2650.stack[3][6] ),
    .B1(\as2650.stack[2][6] ),
    .B2(_3331_),
    .C(_4488_),
    .ZN(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8280_ (.A1(_3437_),
    .A2(_3439_),
    .B1(_3441_),
    .B2(_3442_),
    .ZN(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8281_ (.I(_2210_),
    .Z(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8282_ (.A1(_2241_),
    .A2(_3416_),
    .B1(_3443_),
    .B2(_3444_),
    .ZN(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8283_ (.A1(_3212_),
    .A2(_3445_),
    .ZN(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8284_ (.A1(_3095_),
    .A2(_3416_),
    .B1(_3436_),
    .B2(_3446_),
    .C(_3299_),
    .ZN(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8285_ (.A1(_1105_),
    .A2(_3341_),
    .B(_3447_),
    .C(_3254_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8286_ (.A1(\as2650.pc[6] ),
    .A2(_2593_),
    .A3(_3381_),
    .ZN(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8287_ (.A1(_1112_),
    .A2(_3448_),
    .Z(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8288_ (.I(_3449_),
    .ZN(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8289_ (.A1(_2184_),
    .A2(_2703_),
    .ZN(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8290_ (.A1(_1112_),
    .A2(_2604_),
    .B(_3451_),
    .ZN(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8291_ (.A1(_3224_),
    .A2(_3452_),
    .ZN(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8292_ (.A1(_1544_),
    .A2(_2335_),
    .B1(_2197_),
    .B2(_2187_),
    .ZN(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8293_ (.A1(_2574_),
    .A2(_3450_),
    .B(_3453_),
    .C(_3454_),
    .ZN(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8294_ (.A1(_1104_),
    .A2(_3424_),
    .ZN(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8295_ (.A1(_2689_),
    .A2(_3456_),
    .Z(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8296_ (.A1(_1189_),
    .A2(_3455_),
    .B1(_3457_),
    .B2(_3310_),
    .ZN(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8297_ (.A1(_1596_),
    .A2(_0747_),
    .Z(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8298_ (.A1(_2649_),
    .A2(_0747_),
    .Z(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _8299_ (.A1(_3459_),
    .A2(_3430_),
    .B(_3460_),
    .ZN(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8300_ (.A1(_0901_),
    .A2(_4363_),
    .A3(_3461_),
    .Z(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8301_ (.A1(_2528_),
    .A2(_3462_),
    .ZN(_3463_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8302_ (.A1(_1545_),
    .A2(_2578_),
    .B(_3384_),
    .C(_3463_),
    .ZN(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8303_ (.A1(_3233_),
    .A2(_3450_),
    .B1(_3458_),
    .B2(_3069_),
    .C(_3464_),
    .ZN(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8304_ (.A1(_3092_),
    .A2(_3465_),
    .ZN(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8305_ (.A1(_3138_),
    .A2(_3449_),
    .B1(_3452_),
    .B2(_2586_),
    .C(_2839_),
    .ZN(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8306_ (.A1(_0386_),
    .A2(\as2650.stack[5][7] ),
    .B1(\as2650.stack[4][7] ),
    .B2(_0383_),
    .ZN(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8307_ (.A1(_3327_),
    .A2(_3468_),
    .Z(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _8308_ (.A1(\as2650.stack[6][7] ),
    .A2(_3200_),
    .B1(_3202_),
    .B2(\as2650.stack[7][7] ),
    .C(_0501_),
    .ZN(_3470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8309_ (.A1(_1582_),
    .A2(\as2650.stack[1][7] ),
    .B1(\as2650.stack[0][7] ),
    .B2(_3238_),
    .ZN(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8310_ (.A1(_3196_),
    .A2(_3471_),
    .Z(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _8311_ (.A1(_0918_),
    .A2(\as2650.stack[3][7] ),
    .B1(\as2650.stack[2][7] ),
    .B2(_3200_),
    .C(_3241_),
    .ZN(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _8312_ (.A1(_3469_),
    .A2(_3470_),
    .B1(_3472_),
    .B2(_3473_),
    .ZN(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8313_ (.A1(_3218_),
    .A2(_3449_),
    .B1(_3474_),
    .B2(_3369_),
    .ZN(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8314_ (.A1(_3466_),
    .A2(_3467_),
    .B(_3475_),
    .ZN(_3476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8315_ (.A1(_3343_),
    .A2(_3476_),
    .ZN(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8316_ (.A1(_3255_),
    .A2(_3449_),
    .B(_3166_),
    .ZN(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8317_ (.A1(_1112_),
    .A2(_3341_),
    .B1(_3477_),
    .B2(_3478_),
    .C(_3122_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _8318_ (.A1(_1111_),
    .A2(_3448_),
    .ZN(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8319_ (.A1(_0967_),
    .A2(_3479_),
    .Z(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8320_ (.I(_3480_),
    .Z(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8321_ (.A1(_2689_),
    .A2(_3456_),
    .ZN(_3482_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8322_ (.A1(_0967_),
    .A2(_3482_),
    .ZN(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8323_ (.I0(_3480_),
    .I1(_3483_),
    .S(_2298_),
    .Z(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8324_ (.A1(_2605_),
    .A2(_2767_),
    .ZN(_3485_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8325_ (.A1(_0967_),
    .A2(_2605_),
    .B(_3485_),
    .ZN(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _8326_ (.A1(_2162_),
    .A2(_2677_),
    .B1(_2198_),
    .B2(_1550_),
    .C(_1577_),
    .ZN(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8327_ (.A1(_2315_),
    .A2(_3480_),
    .ZN(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8328_ (.A1(_3085_),
    .A2(_3486_),
    .B(_3487_),
    .C(_3488_),
    .ZN(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8329_ (.A1(_2615_),
    .A2(_3484_),
    .B(_3489_),
    .C(_3064_),
    .ZN(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8330_ (.A1(_0900_),
    .A2(_4363_),
    .ZN(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8331_ (.A1(_0900_),
    .A2(_4363_),
    .ZN(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _8332_ (.A1(_3491_),
    .A2(_3461_),
    .B(_3492_),
    .ZN(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8333_ (.A1(_2528_),
    .A2(_3493_),
    .ZN(_3494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8334_ (.A1(_2735_),
    .A2(_3494_),
    .ZN(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _8335_ (.A1(_2160_),
    .A2(_2475_),
    .A3(_3493_),
    .ZN(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8336_ (.A1(_3495_),
    .A2(_3496_),
    .ZN(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8337_ (.A1(_3274_),
    .A2(_3497_),
    .ZN(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8338_ (.A1(_3274_),
    .A2(_3481_),
    .B(_3498_),
    .C(_3089_),
    .ZN(_3499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8339_ (.A1(_2991_),
    .A2(_3486_),
    .ZN(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8340_ (.A1(_3097_),
    .A2(_3481_),
    .B(_3500_),
    .C(_3092_),
    .ZN(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8341_ (.A1(_3063_),
    .A2(_3490_),
    .A3(_3499_),
    .A4(_3501_),
    .ZN(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8342_ (.I(_2241_),
    .Z(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8343_ (.A1(_4501_),
    .A2(_3444_),
    .B1(_3503_),
    .B2(_3481_),
    .ZN(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8344_ (.A1(_2940_),
    .A2(_3504_),
    .ZN(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8345_ (.A1(_3255_),
    .A2(_3481_),
    .B1(_3502_),
    .B2(_3505_),
    .C(_3300_),
    .ZN(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8346_ (.A1(_0968_),
    .A2(_3303_),
    .B(_3033_),
    .ZN(_3507_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8347_ (.A1(_3506_),
    .A2(_3507_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _8348_ (.A1(\as2650.pc[9] ),
    .A2(\as2650.pc[8] ),
    .A3(_3479_),
    .ZN(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8349_ (.A1(_0966_),
    .A2(_3479_),
    .ZN(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8350_ (.A1(_0986_),
    .A2(_3509_),
    .ZN(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8351_ (.A1(_3508_),
    .A2(_3510_),
    .ZN(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8352_ (.I(_3511_),
    .Z(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8353_ (.A1(_2803_),
    .A2(_3496_),
    .Z(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8354_ (.A1(_3066_),
    .A2(_3513_),
    .ZN(_3514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8355_ (.A1(_3066_),
    .A2(_3512_),
    .B(_3514_),
    .C(_3183_),
    .ZN(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8356_ (.A1(_0966_),
    .A2(_1110_),
    .A3(_3456_),
    .ZN(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8357_ (.A1(_0986_),
    .A2(_3516_),
    .Z(_3517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8358_ (.A1(_3263_),
    .A2(_3517_),
    .B(_3064_),
    .ZN(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8359_ (.A1(_2315_),
    .A2(_3511_),
    .ZN(_3519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8360_ (.A1(_0986_),
    .A2(_3171_),
    .ZN(_3520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8361_ (.A1(_1621_),
    .A2(_2792_),
    .B(_3520_),
    .ZN(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8362_ (.A1(_2784_),
    .A2(_3222_),
    .B1(_3521_),
    .B2(_3419_),
    .ZN(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8363_ (.A1(_3519_),
    .A2(_3522_),
    .B(_3010_),
    .ZN(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8364_ (.A1(_3038_),
    .A2(_3512_),
    .B(_3518_),
    .C(_3523_),
    .ZN(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8365_ (.A1(_3138_),
    .A2(_3512_),
    .B1(_3521_),
    .B2(_2573_),
    .C(_2838_),
    .ZN(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8366_ (.A1(_0398_),
    .A2(_3100_),
    .B1(_3077_),
    .B2(_3511_),
    .C(_2939_),
    .ZN(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _8367_ (.A1(_3515_),
    .A2(_3524_),
    .A3(_3525_),
    .B(_3526_),
    .ZN(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8368_ (.I(_3302_),
    .Z(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8369_ (.A1(_3343_),
    .A2(_3512_),
    .B(_3527_),
    .C(_3528_),
    .ZN(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8370_ (.A1(_2777_),
    .A2(_3303_),
    .B(_3529_),
    .ZN(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8371_ (.A1(_3123_),
    .A2(_3530_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8372_ (.A1(_0998_),
    .A2(_3508_),
    .Z(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8373_ (.I(_3531_),
    .Z(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8374_ (.A1(_0985_),
    .A2(_3516_),
    .ZN(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8375_ (.A1(_2815_),
    .A2(_3533_),
    .Z(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _8376_ (.A1(_3089_),
    .A2(_3263_),
    .A3(_3534_),
    .B(_3034_),
    .ZN(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8377_ (.A1(_2217_),
    .A2(_2934_),
    .ZN(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8378_ (.A1(_2803_),
    .A2(_3496_),
    .ZN(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8379_ (.A1(_2168_),
    .A2(_3537_),
    .ZN(_3538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8380_ (.A1(_2814_),
    .A2(_2320_),
    .ZN(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8381_ (.A1(_2426_),
    .A2(_2846_),
    .B(_3539_),
    .ZN(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8382_ (.A1(_2168_),
    .A2(_2236_),
    .ZN(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8383_ (.A1(_3281_),
    .A2(_3541_),
    .B(_2601_),
    .ZN(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8384_ (.A1(_3419_),
    .A2(_3540_),
    .B1(_3531_),
    .B2(_2961_),
    .C(_3542_),
    .ZN(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8385_ (.A1(_3536_),
    .A2(_3538_),
    .B1(_3543_),
    .B2(_3183_),
    .ZN(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8386_ (.A1(_3347_),
    .A2(_3532_),
    .B1(_3544_),
    .B2(_1639_),
    .ZN(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8387_ (.A1(_2348_),
    .A2(_3540_),
    .B1(_3532_),
    .B2(_3128_),
    .C(_3191_),
    .ZN(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8388_ (.A1(_3535_),
    .A2(_3545_),
    .B(_3546_),
    .ZN(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8389_ (.I(_3532_),
    .ZN(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8390_ (.A1(_0505_),
    .A2(_3369_),
    .B1(_3287_),
    .B2(_3548_),
    .C(_3251_),
    .ZN(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8391_ (.A1(_3095_),
    .A2(_3532_),
    .B1(_3547_),
    .B2(_3549_),
    .C(_3299_),
    .ZN(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8392_ (.I(_1693_),
    .Z(_3551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8393_ (.I(_3551_),
    .Z(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8394_ (.A1(_0998_),
    .A2(_3341_),
    .B(_3550_),
    .C(_3552_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _8395_ (.A1(_0997_),
    .A2(_3508_),
    .ZN(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8396_ (.A1(_2855_),
    .A2(_3553_),
    .Z(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8397_ (.I(_3554_),
    .Z(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8398_ (.A1(_2169_),
    .A2(_3537_),
    .ZN(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8399_ (.A1(_2173_),
    .A2(_3556_),
    .Z(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8400_ (.I0(_2855_),
    .I1(_2879_),
    .S(_2604_),
    .Z(_3558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8401_ (.A1(_2172_),
    .A2(_2778_),
    .ZN(_3559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8402_ (.A1(_3559_),
    .A2(_3322_),
    .B(_2217_),
    .ZN(_3560_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8403_ (.A1(_2315_),
    .A2(_3554_),
    .B1(_3558_),
    .B2(_3419_),
    .C(_3560_),
    .ZN(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8404_ (.A1(_3536_),
    .A2(_3557_),
    .B1(_3561_),
    .B2(_2935_),
    .ZN(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8405_ (.A1(_3347_),
    .A2(_3555_),
    .B1(_3562_),
    .B2(_1639_),
    .ZN(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8406_ (.A1(_2839_),
    .A2(_3563_),
    .ZN(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8407_ (.A1(_2531_),
    .A2(_3558_),
    .ZN(_3565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8408_ (.A1(_1395_),
    .A2(_3555_),
    .ZN(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8409_ (.A1(_3091_),
    .A2(_3565_),
    .A3(_3566_),
    .ZN(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8410_ (.A1(_2815_),
    .A2(_3533_),
    .ZN(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8411_ (.A1(_2856_),
    .A2(_3568_),
    .Z(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8412_ (.A1(_3064_),
    .A2(_3310_),
    .A3(_3569_),
    .ZN(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8413_ (.A1(_3567_),
    .A2(_3570_),
    .ZN(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8414_ (.A1(_3503_),
    .A2(_3555_),
    .B(_3342_),
    .ZN(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8415_ (.A1(_0597_),
    .A2(_3101_),
    .B1(_3571_),
    .B2(_3114_),
    .C(_3572_),
    .ZN(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8416_ (.A1(_3255_),
    .A2(_3555_),
    .B1(_3564_),
    .B2(_3573_),
    .C(_3300_),
    .ZN(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8417_ (.A1(_2856_),
    .A2(_3303_),
    .B(_3033_),
    .ZN(_3575_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8418_ (.A1(_3574_),
    .A2(_3575_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8419_ (.A1(_2854_),
    .A2(_3553_),
    .ZN(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8420_ (.A1(_1017_),
    .A2(_3576_),
    .Z(_3577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8421_ (.I(_3577_),
    .Z(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8422_ (.A1(_2855_),
    .A2(_2814_),
    .A3(_3533_),
    .ZN(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8423_ (.A1(_1018_),
    .A2(_3579_),
    .Z(_3580_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8424_ (.A1(\as2650.addr_buff[3] ),
    .A2(_2333_),
    .A3(_2820_),
    .A4(_3493_),
    .ZN(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8425_ (.A1(_2903_),
    .A2(_3581_),
    .Z(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8426_ (.A1(_2144_),
    .A2(_3582_),
    .ZN(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8427_ (.A1(_2886_),
    .A2(_1543_),
    .ZN(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8428_ (.A1(_1616_),
    .A2(_2910_),
    .B(_3584_),
    .ZN(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8429_ (.A1(_2177_),
    .A2(_2334_),
    .B(_3349_),
    .ZN(_3586_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8430_ (.A1(_2216_),
    .A2(_3586_),
    .B(_2150_),
    .ZN(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8431_ (.A1(_3357_),
    .A2(_3577_),
    .B1(_3585_),
    .B2(_3224_),
    .C(_3587_),
    .ZN(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8432_ (.A1(_3583_),
    .A2(_3588_),
    .ZN(_3589_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _8433_ (.A1(_3088_),
    .A2(_3231_),
    .A3(_3580_),
    .B1(_3589_),
    .B2(_1638_),
    .ZN(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8434_ (.A1(_3137_),
    .A2(_3578_),
    .B1(_3585_),
    .B2(_2572_),
    .C(_2837_),
    .ZN(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8435_ (.A1(_2970_),
    .A2(_3590_),
    .B(_3591_),
    .ZN(_3592_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8436_ (.A1(_3347_),
    .A2(_3578_),
    .B1(_3592_),
    .B2(_2245_),
    .ZN(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8437_ (.A1(_0708_),
    .A2(_3369_),
    .ZN(_3594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8438_ (.A1(_3593_),
    .A2(_3594_),
    .ZN(_3595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8439_ (.A1(_3343_),
    .A2(_3578_),
    .B(_3595_),
    .ZN(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8440_ (.A1(_3078_),
    .A2(_3578_),
    .B(_3166_),
    .ZN(_3597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8441_ (.A1(_1018_),
    .A2(_3300_),
    .B1(_3596_),
    .B2(_3597_),
    .C(_3122_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8442_ (.I(_0781_),
    .ZN(_3598_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8443_ (.A1(_2886_),
    .A2(_2854_),
    .A3(_3553_),
    .ZN(_3599_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8444_ (.A1(\as2650.pc[13] ),
    .A2(_3599_),
    .ZN(_3600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8445_ (.I(_3600_),
    .Z(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8446_ (.A1(_2903_),
    .A2(_3581_),
    .B(_3396_),
    .C(_3273_),
    .ZN(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8447_ (.A1(_2841_),
    .A2(_3601_),
    .B(_3602_),
    .ZN(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8448_ (.A1(\as2650.pc[13] ),
    .A2(_1620_),
    .Z(_3604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8449_ (.A1(_3138_),
    .A2(_3600_),
    .B1(_3604_),
    .B2(_2572_),
    .C(_2838_),
    .ZN(_3605_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8450_ (.A1(_1018_),
    .A2(_3579_),
    .ZN(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8451_ (.A1(_1025_),
    .A2(_3606_),
    .Z(_3607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8452_ (.A1(_3357_),
    .A2(_3600_),
    .ZN(_3608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8453_ (.A1(_2180_),
    .A2(_2335_),
    .B1(_3360_),
    .B2(_3604_),
    .C(_2960_),
    .ZN(_3609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8454_ (.A1(_3608_),
    .A2(_3609_),
    .ZN(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8455_ (.A1(_3266_),
    .A2(_3601_),
    .B1(_3607_),
    .B2(_3310_),
    .C(_3610_),
    .ZN(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8456_ (.A1(_3069_),
    .A2(_3603_),
    .B(_3605_),
    .C(_3611_),
    .ZN(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8457_ (.A1(_3598_),
    .A2(_3101_),
    .B1(_3287_),
    .B2(_3601_),
    .C(_3612_),
    .ZN(_3613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8458_ (.A1(_3212_),
    .A2(_3601_),
    .ZN(_3614_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8459_ (.A1(_3095_),
    .A2(_3613_),
    .B(_3614_),
    .C(_3528_),
    .ZN(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8460_ (.A1(_1025_),
    .A2(_3528_),
    .B(_3615_),
    .ZN(_3616_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8461_ (.A1(_3123_),
    .A2(_3616_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8462_ (.A1(\as2650.pc[13] ),
    .A2(\as2650.pc[12] ),
    .A3(_2854_),
    .A4(_3553_),
    .ZN(_3617_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8463_ (.A1(\as2650.pc[14] ),
    .A2(_3617_),
    .ZN(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8464_ (.I(_3618_),
    .Z(_3619_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8465_ (.I(_3619_),
    .ZN(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8466_ (.A1(_1030_),
    .A2(_2768_),
    .A3(_2573_),
    .ZN(_3621_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8467_ (.A1(_3128_),
    .A2(_3620_),
    .B(_3621_),
    .C(_3191_),
    .ZN(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8468_ (.A1(_1025_),
    .A2(_3606_),
    .ZN(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8469_ (.A1(_1030_),
    .A2(_3623_),
    .ZN(_3624_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8470_ (.A1(\as2650.pc[14] ),
    .A2(_1620_),
    .A3(_2420_),
    .ZN(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8471_ (.A1(_1350_),
    .A2(_3625_),
    .ZN(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8472_ (.A1(_2182_),
    .A2(_2335_),
    .B1(_3357_),
    .B2(_3618_),
    .C(_3626_),
    .ZN(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8473_ (.A1(_3266_),
    .A2(_3620_),
    .B(_3627_),
    .C(_2960_),
    .ZN(_3628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8474_ (.A1(_3263_),
    .A2(_3624_),
    .B(_3628_),
    .ZN(_3629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8475_ (.A1(_2841_),
    .A2(_3421_),
    .ZN(_3630_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8476_ (.A1(_3274_),
    .A2(_3619_),
    .B(_3630_),
    .C(_2960_),
    .ZN(_3631_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8477_ (.A1(_3034_),
    .A2(_3629_),
    .A3(_3631_),
    .ZN(_3632_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8478_ (.A1(_0854_),
    .A2(_3444_),
    .ZN(_3633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8479_ (.A1(_3287_),
    .A2(_3619_),
    .B1(_3622_),
    .B2(_3632_),
    .C(_3633_),
    .ZN(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8480_ (.A1(_3212_),
    .A2(_3619_),
    .ZN(_3635_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8481_ (.A1(_2940_),
    .A2(_3634_),
    .B(_3635_),
    .C(_3302_),
    .ZN(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8482_ (.A1(_1030_),
    .A2(_3528_),
    .B(_3636_),
    .ZN(_3637_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8483_ (.A1(_3123_),
    .A2(_3637_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8484_ (.I(_2436_),
    .Z(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8485_ (.I(_2779_),
    .Z(_3639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8486_ (.I(_2207_),
    .Z(_3640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8487_ (.I(_3640_),
    .Z(_3641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8488_ (.A1(_2362_),
    .A2(_4438_),
    .ZN(_3642_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8489_ (.A1(_3139_),
    .A2(_4459_),
    .B(_2370_),
    .C(_3642_),
    .ZN(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8490_ (.A1(_3639_),
    .A2(_4347_),
    .B1(_3641_),
    .B2(_3643_),
    .ZN(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8491_ (.A1(_1187_),
    .A2(_3209_),
    .ZN(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8492_ (.I(_4152_),
    .Z(_3646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8493_ (.I(_3646_),
    .Z(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8494_ (.I(_2273_),
    .Z(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8495_ (.A1(_4478_),
    .A2(_2956_),
    .ZN(_3649_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8496_ (.A1(_4335_),
    .A2(_3648_),
    .B(_3649_),
    .ZN(_3650_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8497_ (.A1(_3647_),
    .A2(_0962_),
    .B1(_3650_),
    .B2(_4169_),
    .ZN(_3651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8498_ (.I(_1519_),
    .Z(_3652_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8499_ (.A1(_3645_),
    .A2(_3651_),
    .B(_3652_),
    .ZN(_3653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8500_ (.A1(_1516_),
    .A2(_3653_),
    .B(_1535_),
    .ZN(_3654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8501_ (.A1(_1538_),
    .A2(_0441_),
    .B(_3654_),
    .C(_1546_),
    .ZN(_3655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8502_ (.A1(_1669_),
    .A2(_1548_),
    .B(_3655_),
    .C(_3062_),
    .ZN(_3656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8503_ (.A1(_3063_),
    .A2(_4399_),
    .B(_3656_),
    .C(_1632_),
    .ZN(_3657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _8504_ (.A1(_2280_),
    .A2(_2497_),
    .B(_2288_),
    .ZN(_3658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _8505_ (.A1(_1485_),
    .A2(_2125_),
    .B(_2923_),
    .C(_4265_),
    .ZN(_3659_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _8506_ (.A1(_0333_),
    .A2(_4392_),
    .A3(_4514_),
    .A4(_1362_),
    .ZN(_3660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8507_ (.A1(_1435_),
    .A2(_2202_),
    .B(_1468_),
    .C(_1380_),
    .ZN(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8508_ (.A1(_3646_),
    .A2(_1576_),
    .A3(_3660_),
    .A4(_3661_),
    .ZN(_3662_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8509_ (.A1(_4243_),
    .A2(_4244_),
    .A3(_4426_),
    .ZN(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8510_ (.A1(_2333_),
    .A2(_4263_),
    .B1(_4424_),
    .B2(_3663_),
    .ZN(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8511_ (.A1(_4251_),
    .A2(_3664_),
    .ZN(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8512_ (.A1(_1472_),
    .A2(_2261_),
    .B(_3665_),
    .C(_1462_),
    .ZN(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _8513_ (.A1(_0924_),
    .A2(_1449_),
    .A3(_2235_),
    .A4(_1444_),
    .ZN(_3667_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _8514_ (.A1(_1438_),
    .A2(_3662_),
    .A3(_3666_),
    .A4(_3667_),
    .Z(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8515_ (.A1(_1033_),
    .A2(_2155_),
    .A3(_3659_),
    .A4(_3668_),
    .ZN(_3669_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _8516_ (.A1(_1511_),
    .A2(_4405_),
    .A3(_4269_),
    .A4(_2279_),
    .Z(_3670_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8517_ (.A1(_4269_),
    .A2(_4248_),
    .B(_4234_),
    .ZN(_3671_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8518_ (.A1(_1154_),
    .A2(_1433_),
    .B(_3671_),
    .C(_4203_),
    .ZN(_3672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8519_ (.A1(_1197_),
    .A2(_3672_),
    .ZN(_3673_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8520_ (.A1(_1252_),
    .A2(_4278_),
    .A3(_1453_),
    .ZN(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _8521_ (.A1(_4141_),
    .A2(_1197_),
    .A3(_0969_),
    .B(_2148_),
    .ZN(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8522_ (.A1(_3670_),
    .A2(_3673_),
    .A3(_3674_),
    .A4(_3675_),
    .ZN(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _8523_ (.A1(_2265_),
    .A2(_3658_),
    .A3(_3669_),
    .A4(_3676_),
    .ZN(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8524_ (.I(_3677_),
    .Z(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8525_ (.A1(_0368_),
    .A2(_2373_),
    .B(_3678_),
    .ZN(_3679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8526_ (.I(_3677_),
    .Z(_3680_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _8527_ (.A1(_3644_),
    .A2(_3657_),
    .A3(_3679_),
    .B1(_3680_),
    .B2(_1054_),
    .ZN(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8528_ (.A1(_3638_),
    .A2(_3681_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8529_ (.I(_3677_),
    .ZN(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8530_ (.I(_3682_),
    .Z(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8531_ (.I(_1564_),
    .Z(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8532_ (.A1(_2983_),
    .A2(_0328_),
    .Z(_3685_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8533_ (.A1(_3139_),
    .A2(_0320_),
    .B(_2439_),
    .C(_3685_),
    .ZN(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8534_ (.A1(_3639_),
    .A2(_0313_),
    .B1(_3640_),
    .B2(_3686_),
    .ZN(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8535_ (.I(_1514_),
    .Z(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8536_ (.I(_1396_),
    .Z(_3689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8537_ (.I(_0348_),
    .Z(_3690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8538_ (.A1(_3646_),
    .A2(_0984_),
    .B(_1519_),
    .ZN(_3691_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8539_ (.A1(_1492_),
    .A2(_2956_),
    .ZN(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8540_ (.A1(_3328_),
    .A2(_2956_),
    .B(_3692_),
    .C(_4507_),
    .ZN(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8541_ (.A1(_4507_),
    .A2(_3249_),
    .B(_3693_),
    .C(_1376_),
    .ZN(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8542_ (.A1(_3652_),
    .A2(_0367_),
    .B1(_3691_),
    .B2(_3694_),
    .ZN(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8543_ (.A1(_3689_),
    .A2(_3695_),
    .ZN(_3696_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8544_ (.A1(_3689_),
    .A2(_3690_),
    .B(_3696_),
    .C(_1514_),
    .ZN(_3697_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8545_ (.A1(_1680_),
    .A2(_3688_),
    .B(_3697_),
    .C(_2411_),
    .ZN(_3698_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8546_ (.A1(_0361_),
    .A2(_1677_),
    .B(_3678_),
    .C(_3698_),
    .ZN(_3699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8547_ (.A1(_1200_),
    .A2(_3684_),
    .B(_3687_),
    .C(_3699_),
    .ZN(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8548_ (.A1(_3003_),
    .A2(_3683_),
    .B(_3700_),
    .C(_3552_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8549_ (.I(_2983_),
    .Z(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8550_ (.A1(_2648_),
    .A2(_0485_),
    .ZN(_3702_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8551_ (.A1(_3701_),
    .A2(_0476_),
    .B(_2557_),
    .C(_3702_),
    .ZN(_3703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8552_ (.A1(_3639_),
    .A2(_0437_),
    .B1(_3641_),
    .B2(_3703_),
    .ZN(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8553_ (.I(_3646_),
    .Z(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8554_ (.A1(\as2650.overflow ),
    .A2(_3648_),
    .ZN(_3706_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8555_ (.A1(_1400_),
    .A2(_1348_),
    .A3(_1403_),
    .ZN(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8556_ (.A1(\as2650.psu[2] ),
    .A2(_3707_),
    .B(_4465_),
    .ZN(_3708_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8557_ (.A1(_1187_),
    .A2(_3297_),
    .B1(_3706_),
    .B2(_3708_),
    .C(_3647_),
    .ZN(_3709_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8558_ (.A1(_3705_),
    .A2(_0996_),
    .B(_3709_),
    .C(_3652_),
    .ZN(_3710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8559_ (.A1(_1517_),
    .A2(_1200_),
    .ZN(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8560_ (.A1(_3710_),
    .A2(_3711_),
    .B(_1535_),
    .ZN(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8561_ (.I(_1396_),
    .Z(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8562_ (.A1(_3713_),
    .A2(_0681_),
    .B(_1515_),
    .ZN(_3714_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8563_ (.A1(_1683_),
    .A2(_3688_),
    .B1(_3712_),
    .B2(_3714_),
    .C(_2411_),
    .ZN(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8564_ (.A1(_3690_),
    .A2(_2373_),
    .B1(_2533_),
    .B2(_0463_),
    .C(_3715_),
    .ZN(_3716_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8565_ (.A1(_3682_),
    .A2(_3704_),
    .A3(_3716_),
    .ZN(_3717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8566_ (.A1(_1254_),
    .A2(_3683_),
    .B(_3717_),
    .C(_3552_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8567_ (.I(_3689_),
    .Z(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8568_ (.I(_4409_),
    .Z(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8569_ (.I(_2273_),
    .Z(_3720_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8570_ (.A1(_4357_),
    .A2(_3720_),
    .ZN(_3721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8571_ (.I(_4506_),
    .Z(_3722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8572_ (.A1(_1588_),
    .A2(_2957_),
    .B(_3721_),
    .C(_3722_),
    .ZN(_3723_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8573_ (.I(_1376_),
    .Z(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8574_ (.A1(_4508_),
    .A2(_3337_),
    .B(_3723_),
    .C(_3724_),
    .ZN(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8575_ (.A1(_3705_),
    .A2(_1007_),
    .B(_3719_),
    .ZN(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8576_ (.A1(_3719_),
    .A2(_3690_),
    .B1(_3725_),
    .B2(_3726_),
    .C(_3713_),
    .ZN(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8577_ (.A1(_3718_),
    .A2(_0742_),
    .B(_3727_),
    .C(_1574_),
    .ZN(_3728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8578_ (.A1(_2171_),
    .A2(_1548_),
    .ZN(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8579_ (.A1(_3728_),
    .A2(_3729_),
    .ZN(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8580_ (.A1(_0681_),
    .A2(_1446_),
    .B1(_2533_),
    .B2(_0560_),
    .C(_3677_),
    .ZN(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8581_ (.A1(_2648_),
    .A2(_0580_),
    .ZN(_3732_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8582_ (.A1(_3701_),
    .A2(_0575_),
    .B(_2557_),
    .C(_3732_),
    .ZN(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8583_ (.A1(_3639_),
    .A2(_0541_),
    .B1(_3641_),
    .B2(_3733_),
    .ZN(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8584_ (.A1(_2239_),
    .A2(_3730_),
    .B(_3731_),
    .C(_3734_),
    .ZN(_3735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8585_ (.A1(_3014_),
    .A2(_3683_),
    .B(_3735_),
    .C(_3552_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8586_ (.A1(_2983_),
    .A2(_0686_),
    .Z(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8587_ (.A1(_2362_),
    .A2(_0643_),
    .B(_2439_),
    .C(_3736_),
    .ZN(_3737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8588_ (.A1(_2779_),
    .A2(_0634_),
    .B1(_3640_),
    .B2(_3737_),
    .ZN(_3738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8589_ (.A1(_0673_),
    .A2(_2797_),
    .ZN(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8590_ (.A1(_1229_),
    .A2(_2957_),
    .ZN(_3740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8591_ (.A1(\as2650.psu[4] ),
    .A2(_3707_),
    .B(_4465_),
    .ZN(_3741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8592_ (.A1(_3722_),
    .A2(_3376_),
    .ZN(_3742_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8593_ (.A1(_3740_),
    .A2(_3741_),
    .B(_3647_),
    .C(_3742_),
    .ZN(_3743_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8594_ (.A1(_3705_),
    .A2(_1016_),
    .B(_3743_),
    .C(_1520_),
    .ZN(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8595_ (.A1(_1517_),
    .A2(_0557_),
    .ZN(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8596_ (.A1(_3744_),
    .A2(_3745_),
    .B(_1538_),
    .ZN(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8597_ (.I(_0665_),
    .Z(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8598_ (.A1(_1575_),
    .A2(_3747_),
    .B(_1515_),
    .ZN(_3748_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8599_ (.A1(_2176_),
    .A2(_3688_),
    .B1(_3746_),
    .B2(_3748_),
    .C(_2411_),
    .ZN(_3749_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8600_ (.A1(_3678_),
    .A2(_3739_),
    .A3(_3749_),
    .ZN(_3750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8601_ (.A1(_0742_),
    .A2(_3684_),
    .B(_3738_),
    .C(_3750_),
    .ZN(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8602_ (.I(_3551_),
    .Z(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8603_ (.A1(_1090_),
    .A2(_3682_),
    .B(_3751_),
    .C(_3752_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8604_ (.A1(_2399_),
    .A2(_0741_),
    .ZN(_3753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8605_ (.A1(_2648_),
    .A2(_0771_),
    .ZN(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8606_ (.A1(_2557_),
    .A2(_3753_),
    .A3(_3754_),
    .ZN(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8607_ (.A1(_2779_),
    .A2(_0736_),
    .B1(_3640_),
    .B2(_3755_),
    .ZN(_3756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8608_ (.A1(_1538_),
    .A2(_0792_),
    .ZN(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8609_ (.A1(\as2650.psu[5] ),
    .A2(_3648_),
    .ZN(_3758_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8610_ (.A1(_1602_),
    .A2(_3720_),
    .B(_3758_),
    .ZN(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8611_ (.A1(_4507_),
    .A2(_3410_),
    .Z(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _8612_ (.A1(_3724_),
    .A2(_1024_),
    .B1(_3759_),
    .B2(_0695_),
    .C(_3760_),
    .ZN(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8613_ (.A1(_1360_),
    .A2(_0638_),
    .ZN(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8614_ (.A1(_1517_),
    .A2(_3761_),
    .B(_3762_),
    .ZN(_3763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8615_ (.A1(_3689_),
    .A2(_3763_),
    .B(_1546_),
    .ZN(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8616_ (.A1(_2179_),
    .A2(_1546_),
    .B1(_3757_),
    .B2(_3764_),
    .C(_3062_),
    .ZN(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8617_ (.A1(_3114_),
    .A2(_2293_),
    .B(_3765_),
    .C(_2772_),
    .ZN(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8618_ (.A1(_3747_),
    .A2(_3684_),
    .B(_3756_),
    .C(_3766_),
    .ZN(_3767_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8619_ (.A1(_3682_),
    .A2(_3767_),
    .B(_2230_),
    .ZN(_3768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8620_ (.A1(_0651_),
    .A2(_3683_),
    .B(_3768_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8621_ (.A1(_2399_),
    .A2(_0841_),
    .Z(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8622_ (.A1(_3701_),
    .A2(_0821_),
    .B(_2385_),
    .C(_3769_),
    .ZN(_3770_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8623_ (.A1(_3079_),
    .A2(_0814_),
    .B1(_2208_),
    .B2(_3770_),
    .ZN(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8624_ (.A1(_3705_),
    .A2(_1040_),
    .B(_3652_),
    .ZN(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8625_ (.A1(_1429_),
    .A2(_3720_),
    .ZN(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8626_ (.A1(_1583_),
    .A2(_2957_),
    .B(_3773_),
    .C(_3722_),
    .ZN(_3774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8627_ (.A1(_4508_),
    .A2(_3443_),
    .B(_3774_),
    .C(_3724_),
    .ZN(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8628_ (.A1(_1520_),
    .A2(_3747_),
    .B1(_3772_),
    .B2(_3775_),
    .C(_3713_),
    .ZN(_3776_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8629_ (.A1(_1575_),
    .A2(_4370_),
    .B(_3776_),
    .C(_3688_),
    .ZN(_3777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8630_ (.A1(_1560_),
    .A2(_1548_),
    .B(_2438_),
    .ZN(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8631_ (.A1(_1539_),
    .A2(_3684_),
    .B1(_3777_),
    .B2(_3778_),
    .ZN(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8632_ (.A1(_0829_),
    .A2(_1677_),
    .B(_3771_),
    .C(_3779_),
    .ZN(_3780_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8633_ (.A1(_1102_),
    .A2(_3680_),
    .ZN(_3781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8634_ (.A1(_3680_),
    .A2(_3780_),
    .B(_3781_),
    .C(_3752_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8635_ (.A1(_0862_),
    .A2(_3680_),
    .ZN(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8636_ (.A1(_3079_),
    .A2(_0884_),
    .Z(_3783_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8637_ (.A1(_3701_),
    .A2(_0894_),
    .ZN(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8638_ (.A1(_3139_),
    .A2(_0891_),
    .B(_2370_),
    .ZN(_3785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8639_ (.A1(_3784_),
    .A2(_3785_),
    .B(_3641_),
    .ZN(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8640_ (.A1(_3722_),
    .A2(_3474_),
    .ZN(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8641_ (.A1(\as2650.psu[7] ),
    .A2(_3648_),
    .ZN(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8642_ (.A1(_1619_),
    .A2(_3720_),
    .B(_3788_),
    .ZN(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8643_ (.A1(_1376_),
    .A2(_2082_),
    .B1(_3789_),
    .B2(_0695_),
    .ZN(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8644_ (.A1(_3787_),
    .A2(_3790_),
    .ZN(_3791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8645_ (.A1(_1576_),
    .A2(_3791_),
    .ZN(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8646_ (.A1(_3713_),
    .A2(_0905_),
    .B(_1518_),
    .C(_3792_),
    .ZN(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8647_ (.I(_1547_),
    .ZN(_3794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8648_ (.A1(_1515_),
    .A2(_3793_),
    .B(_3794_),
    .ZN(_3795_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8649_ (.A1(_1636_),
    .A2(_2373_),
    .B1(_3795_),
    .B2(_2438_),
    .C(_3678_),
    .ZN(_3796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8650_ (.A1(_0898_),
    .A2(_2797_),
    .B1(_3783_),
    .B2(_3786_),
    .C(_3796_),
    .ZN(_3797_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8651_ (.A1(_1644_),
    .A2(_3782_),
    .A3(_3797_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8652_ (.A1(_1889_),
    .A2(_1854_),
    .A3(_1118_),
    .ZN(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8653_ (.I(_3798_),
    .Z(_3799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8654_ (.I(_3798_),
    .Z(_3800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8655_ (.A1(\as2650.stack[6][0] ),
    .A2(_3800_),
    .ZN(_3801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8656_ (.A1(_1888_),
    .A2(_3799_),
    .B(_3801_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8657_ (.A1(\as2650.stack[6][1] ),
    .A2(_3800_),
    .ZN(_3802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8658_ (.A1(_1894_),
    .A2(_3799_),
    .B(_3802_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8659_ (.A1(\as2650.stack[6][2] ),
    .A2(_3800_),
    .ZN(_3803_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8660_ (.A1(_1896_),
    .A2(_3799_),
    .B(_3803_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8661_ (.A1(\as2650.stack[6][3] ),
    .A2(_3800_),
    .ZN(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8662_ (.A1(_1898_),
    .A2(_3799_),
    .B(_3804_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8663_ (.I(_3798_),
    .Z(_3805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8664_ (.I(_3798_),
    .Z(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8665_ (.A1(\as2650.stack[6][4] ),
    .A2(_3806_),
    .ZN(_3807_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8666_ (.A1(_1900_),
    .A2(_3805_),
    .B(_3807_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8667_ (.A1(\as2650.stack[6][5] ),
    .A2(_3806_),
    .ZN(_3808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8668_ (.A1(_1904_),
    .A2(_3805_),
    .B(_3808_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8669_ (.A1(\as2650.stack[6][6] ),
    .A2(_3806_),
    .ZN(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8670_ (.A1(_1906_),
    .A2(_3805_),
    .B(_3809_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8671_ (.A1(\as2650.stack[6][7] ),
    .A2(_3806_),
    .ZN(_3810_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8672_ (.A1(_1908_),
    .A2(_3805_),
    .B(_3810_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8673_ (.I(_0976_),
    .Z(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8674_ (.A1(_4495_),
    .A2(_1050_),
    .ZN(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8675_ (.A1(_0917_),
    .A2(_3812_),
    .ZN(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8676_ (.I(_3813_),
    .Z(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8677_ (.I(_3814_),
    .Z(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8678_ (.I(_3814_),
    .Z(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8679_ (.A1(\as2650.stack[5][8] ),
    .A2(_3816_),
    .ZN(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8680_ (.A1(_3811_),
    .A2(_3815_),
    .B(_3817_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8681_ (.I(_0989_),
    .Z(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8682_ (.I(_3813_),
    .Z(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8683_ (.A1(\as2650.stack[5][9] ),
    .A2(_3819_),
    .ZN(_3820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8684_ (.A1(_3818_),
    .A2(_3815_),
    .B(_3820_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8685_ (.I(_1000_),
    .Z(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8686_ (.A1(\as2650.stack[5][10] ),
    .A2(_3819_),
    .ZN(_3822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8687_ (.A1(_3821_),
    .A2(_3815_),
    .B(_3822_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8688_ (.I(_1011_),
    .Z(_3823_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8689_ (.A1(\as2650.stack[5][11] ),
    .A2(_3819_),
    .ZN(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8690_ (.A1(_3823_),
    .A2(_3815_),
    .B(_3824_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8691_ (.I(_1020_),
    .Z(_3825_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8692_ (.A1(\as2650.stack[5][12] ),
    .A2(_3819_),
    .ZN(_3826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8693_ (.A1(_3825_),
    .A2(_3816_),
    .B(_3826_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8694_ (.I(_1027_),
    .Z(_3827_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8695_ (.A1(\as2650.stack[5][13] ),
    .A2(_3814_),
    .ZN(_3828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8696_ (.A1(_3827_),
    .A2(_3816_),
    .B(_3828_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8697_ (.I(_1042_),
    .Z(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8698_ (.A1(\as2650.stack[5][14] ),
    .A2(_3814_),
    .ZN(_3830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8699_ (.A1(_3829_),
    .A2(_3816_),
    .B(_3830_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8700_ (.A1(_0917_),
    .A2(_1047_),
    .A3(_1117_),
    .ZN(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8701_ (.I(_3831_),
    .Z(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8702_ (.I(_3832_),
    .Z(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8703_ (.I(_3832_),
    .Z(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8704_ (.A1(\as2650.stack[4][8] ),
    .A2(_3834_),
    .ZN(_3835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8705_ (.A1(_3811_),
    .A2(_3833_),
    .B(_3835_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8706_ (.I(_3831_),
    .Z(_3836_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8707_ (.A1(\as2650.stack[4][9] ),
    .A2(_3836_),
    .ZN(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8708_ (.A1(_3818_),
    .A2(_3833_),
    .B(_3837_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8709_ (.A1(\as2650.stack[4][10] ),
    .A2(_3836_),
    .ZN(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8710_ (.A1(_3821_),
    .A2(_3833_),
    .B(_3838_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8711_ (.A1(\as2650.stack[4][11] ),
    .A2(_3836_),
    .ZN(_3839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8712_ (.A1(_3823_),
    .A2(_3833_),
    .B(_3839_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8713_ (.A1(\as2650.stack[4][12] ),
    .A2(_3836_),
    .ZN(_3840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8714_ (.A1(_3825_),
    .A2(_3834_),
    .B(_3840_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8715_ (.A1(\as2650.stack[4][13] ),
    .A2(_3832_),
    .ZN(_3841_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8716_ (.A1(_3827_),
    .A2(_3834_),
    .B(_3841_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8717_ (.A1(\as2650.stack[4][14] ),
    .A2(_3832_),
    .ZN(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8718_ (.A1(_3829_),
    .A2(_3834_),
    .B(_3842_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8719_ (.A1(_0920_),
    .A2(_1049_),
    .ZN(_3843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8720_ (.I(_3843_),
    .Z(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8721_ (.I(_3844_),
    .Z(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8722_ (.I(_3844_),
    .Z(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8723_ (.A1(\as2650.stack[3][8] ),
    .A2(_3846_),
    .ZN(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8724_ (.A1(_3811_),
    .A2(_3845_),
    .B(_3847_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8725_ (.I(_3843_),
    .Z(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8726_ (.A1(\as2650.stack[3][9] ),
    .A2(_3848_),
    .ZN(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8727_ (.A1(_3818_),
    .A2(_3845_),
    .B(_3849_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8728_ (.A1(\as2650.stack[3][10] ),
    .A2(_3848_),
    .ZN(_3850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8729_ (.A1(_3821_),
    .A2(_3845_),
    .B(_3850_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8730_ (.A1(\as2650.stack[3][11] ),
    .A2(_3848_),
    .ZN(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8731_ (.A1(_3823_),
    .A2(_3845_),
    .B(_3851_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8732_ (.A1(\as2650.stack[3][12] ),
    .A2(_3848_),
    .ZN(_3852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8733_ (.A1(_3825_),
    .A2(_3846_),
    .B(_3852_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8734_ (.A1(\as2650.stack[3][13] ),
    .A2(_3844_),
    .ZN(_3853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8735_ (.A1(_3827_),
    .A2(_3846_),
    .B(_3853_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8736_ (.A1(\as2650.stack[3][14] ),
    .A2(_3844_),
    .ZN(_3854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8737_ (.A1(_3829_),
    .A2(_3846_),
    .B(_3854_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8738_ (.A1(_1889_),
    .A2(_1854_),
    .A3(_1051_),
    .ZN(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8739_ (.I(_3855_),
    .Z(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8740_ (.I(_3855_),
    .Z(_3857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8741_ (.A1(\as2650.stack[7][0] ),
    .A2(_3857_),
    .ZN(_3858_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8742_ (.A1(_1888_),
    .A2(_3856_),
    .B(_3858_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8743_ (.A1(\as2650.stack[7][1] ),
    .A2(_3857_),
    .ZN(_3859_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8744_ (.A1(_1894_),
    .A2(_3856_),
    .B(_3859_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8745_ (.A1(\as2650.stack[7][2] ),
    .A2(_3857_),
    .ZN(_3860_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8746_ (.A1(_1896_),
    .A2(_3856_),
    .B(_3860_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8747_ (.A1(\as2650.stack[7][3] ),
    .A2(_3857_),
    .ZN(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8748_ (.A1(_1898_),
    .A2(_3856_),
    .B(_3861_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8749_ (.I(_3855_),
    .Z(_3862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8750_ (.I(_3855_),
    .Z(_3863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8751_ (.A1(\as2650.stack[7][4] ),
    .A2(_3863_),
    .ZN(_3864_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8752_ (.A1(_1900_),
    .A2(_3862_),
    .B(_3864_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8753_ (.A1(\as2650.stack[7][5] ),
    .A2(_3863_),
    .ZN(_3865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8754_ (.A1(_1904_),
    .A2(_3862_),
    .B(_3865_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8755_ (.A1(\as2650.stack[7][6] ),
    .A2(_3863_),
    .ZN(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8756_ (.A1(_1906_),
    .A2(_3862_),
    .B(_3866_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8757_ (.A1(\as2650.stack[7][7] ),
    .A2(_3863_),
    .ZN(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8758_ (.A1(_1908_),
    .A2(_3862_),
    .B(_3867_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8759_ (.A1(_1045_),
    .A2(_3812_),
    .ZN(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8760_ (.I(_3868_),
    .Z(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8761_ (.I(_3869_),
    .Z(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8762_ (.I(_3869_),
    .Z(_3871_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8763_ (.A1(\as2650.stack[7][8] ),
    .A2(_3871_),
    .ZN(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8764_ (.A1(_3811_),
    .A2(_3870_),
    .B(_3872_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8765_ (.I(_3868_),
    .Z(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8766_ (.A1(\as2650.stack[7][9] ),
    .A2(_3873_),
    .ZN(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8767_ (.A1(_3818_),
    .A2(_3870_),
    .B(_3874_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8768_ (.A1(\as2650.stack[7][10] ),
    .A2(_3873_),
    .ZN(_3875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8769_ (.A1(_3821_),
    .A2(_3870_),
    .B(_3875_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8770_ (.A1(\as2650.stack[7][11] ),
    .A2(_3873_),
    .ZN(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8771_ (.A1(_3823_),
    .A2(_3870_),
    .B(_3876_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8772_ (.A1(\as2650.stack[7][12] ),
    .A2(_3873_),
    .ZN(_3877_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8773_ (.A1(_3825_),
    .A2(_3871_),
    .B(_3877_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8774_ (.A1(\as2650.stack[7][13] ),
    .A2(_3869_),
    .ZN(_3878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8775_ (.A1(_3827_),
    .A2(_3871_),
    .B(_3878_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8776_ (.A1(\as2650.stack[7][14] ),
    .A2(_3869_),
    .ZN(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8777_ (.A1(_3829_),
    .A2(_3871_),
    .B(_3879_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _8778_ (.A1(_1229_),
    .A2(_1378_),
    .A3(_1375_),
    .B(_4116_),
    .ZN(_3880_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8779_ (.A1(_1450_),
    .A2(_4179_),
    .A3(_4269_),
    .A4(_4446_),
    .ZN(_3881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8780_ (.A1(_4118_),
    .A2(_1168_),
    .ZN(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8781_ (.A1(_4385_),
    .A2(_3881_),
    .A3(_4413_),
    .A4(_3882_),
    .ZN(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8782_ (.A1(_4257_),
    .A2(_4464_),
    .A3(_0335_),
    .ZN(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _8783_ (.A1(_3883_),
    .A2(_4205_),
    .A3(_4430_),
    .A4(_3884_),
    .ZN(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8784_ (.A1(_1695_),
    .A2(_3885_),
    .Z(_3886_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8785_ (.I(_3886_),
    .ZN(_3887_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8786_ (.A1(_3880_),
    .A2(_3887_),
    .ZN(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8787_ (.I(_3888_),
    .Z(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8788_ (.A1(_0698_),
    .A2(_3888_),
    .ZN(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8789_ (.I(_3890_),
    .Z(_3891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8790_ (.A1(\as2650.r123[1][0] ),
    .A2(_3889_),
    .B1(_3891_),
    .B2(_1701_),
    .ZN(_3892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8791_ (.I(_3887_),
    .Z(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8792_ (.I(_3893_),
    .Z(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8793_ (.A1(_4463_),
    .A2(_3894_),
    .ZN(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8794_ (.A1(_3892_),
    .A2(_3895_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8795_ (.A1(\as2650.r123[1][1] ),
    .A2(_3889_),
    .B1(_3891_),
    .B2(_1711_),
    .ZN(_3896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8796_ (.A1(_0374_),
    .A2(_3894_),
    .ZN(_3897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8797_ (.A1(_3896_),
    .A2(_3897_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8798_ (.I(_3890_),
    .Z(_3898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8799_ (.A1(\as2650.r123[1][2] ),
    .A2(_3889_),
    .B1(_3898_),
    .B2(_1722_),
    .ZN(_3899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8800_ (.A1(_0488_),
    .A2(_3894_),
    .ZN(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8801_ (.A1(_3899_),
    .A2(_3900_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8802_ (.I(_3888_),
    .Z(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8803_ (.A1(\as2650.r123[1][3] ),
    .A2(_3901_),
    .B1(_3898_),
    .B2(_1743_),
    .ZN(_3902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8804_ (.A1(_0583_),
    .A2(_3894_),
    .ZN(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8805_ (.A1(_3902_),
    .A2(_3903_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8806_ (.A1(_3880_),
    .A2(_3887_),
    .B(_4517_),
    .ZN(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8807_ (.A1(_1761_),
    .A2(_3904_),
    .ZN(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8808_ (.A1(\as2650.r123[1][4] ),
    .A2(_3889_),
    .B(_3905_),
    .ZN(_3906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8809_ (.A1(_0690_),
    .A2(_3893_),
    .ZN(_3907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8810_ (.A1(_3906_),
    .A2(_3907_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8811_ (.A1(\as2650.r123[1][5] ),
    .A2(_3901_),
    .B1(_3898_),
    .B2(_1792_),
    .ZN(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8812_ (.A1(_0774_),
    .A2(_3893_),
    .ZN(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8813_ (.A1(_3908_),
    .A2(_3909_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8814_ (.A1(\as2650.r123[1][6] ),
    .A2(_3901_),
    .B1(_3898_),
    .B2(_1822_),
    .ZN(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8815_ (.A1(_0845_),
    .A2(_3893_),
    .ZN(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8816_ (.A1(_3910_),
    .A2(_3911_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8817_ (.A1(_4290_),
    .A2(_0884_),
    .B(_0915_),
    .ZN(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8818_ (.A1(\as2650.r123[1][7] ),
    .A2(_3901_),
    .B1(_3890_),
    .B2(_1852_),
    .ZN(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8819_ (.A1(_3912_),
    .A2(_3886_),
    .B(_3913_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8820_ (.A1(_3885_),
    .A2(_1367_),
    .ZN(_3914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8821_ (.I(_3914_),
    .Z(_3915_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8822_ (.A1(_3880_),
    .A2(_3914_),
    .ZN(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8823_ (.I(_3916_),
    .Z(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8824_ (.A1(_4463_),
    .A2(_3915_),
    .B1(_3917_),
    .B2(\as2650.r123[2][0] ),
    .ZN(_3918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8825_ (.I(_3890_),
    .Z(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8826_ (.A1(_1953_),
    .A2(_3919_),
    .ZN(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8827_ (.A1(_3918_),
    .A2(_3920_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8828_ (.A1(_0374_),
    .A2(_3915_),
    .B1(_3917_),
    .B2(\as2650.r123[2][1] ),
    .ZN(_3921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8829_ (.A1(_1989_),
    .A2(_3919_),
    .ZN(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8830_ (.A1(_3921_),
    .A2(_3922_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8831_ (.A1(_0488_),
    .A2(_3915_),
    .B1(_3917_),
    .B2(\as2650.r123[2][2] ),
    .ZN(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8832_ (.A1(_2021_),
    .A2(_3919_),
    .ZN(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8833_ (.A1(_3923_),
    .A2(_3924_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8834_ (.A1(_0583_),
    .A2(_3915_),
    .B1(_3917_),
    .B2(\as2650.r123[2][3] ),
    .ZN(_3925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8835_ (.A1(_2049_),
    .A2(_3919_),
    .ZN(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8836_ (.A1(_3925_),
    .A2(_3926_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8837_ (.I(_3914_),
    .Z(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8838_ (.I(_3916_),
    .Z(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8839_ (.A1(_0690_),
    .A2(_3927_),
    .B1(_3928_),
    .B2(\as2650.r123[2][4] ),
    .ZN(_3929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8840_ (.A1(_2071_),
    .A2(_3904_),
    .B(_3929_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8841_ (.A1(_0774_),
    .A2(_3927_),
    .B1(_3928_),
    .B2(\as2650.r123[2][5] ),
    .ZN(_3930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8842_ (.A1(_2091_),
    .A2(_3891_),
    .ZN(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8843_ (.A1(_3930_),
    .A2(_3931_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8844_ (.A1(_0845_),
    .A2(_3927_),
    .B1(_3928_),
    .B2(\as2650.r123[2][6] ),
    .ZN(_3932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8845_ (.A1(_2100_),
    .A2(_3891_),
    .ZN(_3933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8846_ (.A1(_3932_),
    .A2(_3933_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8847_ (.I(_3927_),
    .ZN(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8848_ (.A1(\as2650.r123[2][7] ),
    .A2(_3928_),
    .ZN(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8849_ (.A1(_2105_),
    .A2(_3904_),
    .B1(_3934_),
    .B2(_3912_),
    .C(_3935_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8850_ (.A1(_1512_),
    .A2(_4408_),
    .B1(_1415_),
    .B2(_1436_),
    .ZN(_3936_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _8851_ (.A1(_2154_),
    .A2(_2923_),
    .A3(_3658_),
    .A4(_3936_),
    .ZN(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _8852_ (.A1(_2213_),
    .A2(_2920_),
    .A3(_3670_),
    .A4(_3937_),
    .Z(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8853_ (.I(_3938_),
    .Z(_3939_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8854_ (.A1(_1572_),
    .A2(_4245_),
    .Z(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8855_ (.I(_3940_),
    .Z(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8856_ (.I(_3940_),
    .Z(_3942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8857_ (.A1(_0368_),
    .A2(_3942_),
    .ZN(_3943_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8858_ (.A1(_1054_),
    .A2(_3941_),
    .B(_3943_),
    .ZN(_3944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8859_ (.I(_3938_),
    .Z(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8860_ (.A1(net41),
    .A2(_3945_),
    .ZN(_3946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8861_ (.A1(_3939_),
    .A2(_3944_),
    .B(_3946_),
    .C(_3752_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8862_ (.A1(_0441_),
    .A2(_3942_),
    .ZN(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8863_ (.A1(_1065_),
    .A2(_3941_),
    .B(_3947_),
    .ZN(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8864_ (.A1(net42),
    .A2(_3945_),
    .ZN(_3949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8865_ (.A1(_3939_),
    .A2(_3948_),
    .B(_3949_),
    .C(_3752_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8866_ (.A1(_3690_),
    .A2(_3942_),
    .ZN(_3950_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8867_ (.A1(_0506_),
    .A2(_3941_),
    .B(_3950_),
    .ZN(_3951_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8868_ (.A1(net43),
    .A2(_3945_),
    .ZN(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8869_ (.I(_3551_),
    .Z(_3953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8870_ (.A1(_3939_),
    .A2(_3951_),
    .B(_3952_),
    .C(_3953_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8871_ (.A1(_0681_),
    .A2(_3942_),
    .ZN(_3954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8872_ (.A1(_0598_),
    .A2(_3941_),
    .B(_3954_),
    .ZN(_3955_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8873_ (.A1(net44),
    .A2(_3945_),
    .ZN(_3956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8874_ (.A1(_3939_),
    .A2(_3955_),
    .B(_3956_),
    .C(_3953_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8875_ (.I(_3938_),
    .Z(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8876_ (.I(_3940_),
    .Z(_3958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8877_ (.I(_3940_),
    .Z(_3959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8878_ (.A1(_0553_),
    .A2(_3959_),
    .ZN(_3960_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8879_ (.A1(_0699_),
    .A2(_3958_),
    .B(_3960_),
    .ZN(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8880_ (.I(_3938_),
    .Z(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8881_ (.A1(net45),
    .A2(_3962_),
    .ZN(_3963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8882_ (.A1(_3957_),
    .A2(_3961_),
    .B(_3963_),
    .C(_3953_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8883_ (.A1(_3747_),
    .A2(_3959_),
    .ZN(_3964_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8884_ (.A1(_0784_),
    .A2(_3958_),
    .B(_3964_),
    .ZN(_3965_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8885_ (.A1(net19),
    .A2(_3962_),
    .ZN(_3966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8886_ (.A1(_3957_),
    .A2(_3965_),
    .B(_3966_),
    .C(_3953_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8887_ (.A1(_1539_),
    .A2(_3959_),
    .ZN(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8888_ (.A1(_1102_),
    .A2(_3958_),
    .B(_3967_),
    .ZN(_3968_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8889_ (.A1(net20),
    .A2(_3962_),
    .ZN(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8890_ (.I(_3551_),
    .Z(_3970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8891_ (.A1(_3957_),
    .A2(_3968_),
    .B(_3969_),
    .C(_3970_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8892_ (.A1(_1636_),
    .A2(_3959_),
    .ZN(_3971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8893_ (.A1(_0862_),
    .A2(_3958_),
    .B(_3971_),
    .ZN(_3972_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8894_ (.A1(net21),
    .A2(_3962_),
    .ZN(_3973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8895_ (.A1(_3957_),
    .A2(_3972_),
    .B(_3973_),
    .C(_3970_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8896_ (.A1(_1889_),
    .A2(_1048_),
    .A3(_1118_),
    .ZN(_3974_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8897_ (.I(_3974_),
    .Z(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8898_ (.I(_3974_),
    .Z(_3976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8899_ (.A1(\as2650.stack[2][0] ),
    .A2(_3976_),
    .ZN(_3977_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8900_ (.A1(_3975_),
    .A2(_1062_),
    .B(_3977_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8901_ (.A1(\as2650.stack[2][1] ),
    .A2(_3976_),
    .ZN(_3978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8902_ (.A1(_3975_),
    .A2(_1071_),
    .B(_3978_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8903_ (.A1(\as2650.stack[2][2] ),
    .A2(_3976_),
    .ZN(_3979_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8904_ (.A1(_3975_),
    .A2(_1079_),
    .B(_3979_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8905_ (.A1(\as2650.stack[2][3] ),
    .A2(_3976_),
    .ZN(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8906_ (.A1(_3975_),
    .A2(_1087_),
    .B(_3980_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8907_ (.I(_3974_),
    .Z(_3981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8908_ (.I(_3974_),
    .Z(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8909_ (.A1(\as2650.stack[2][4] ),
    .A2(_3982_),
    .ZN(_3983_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8910_ (.A1(_3981_),
    .A2(_1093_),
    .B(_3983_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8911_ (.A1(\as2650.stack[2][5] ),
    .A2(_3982_),
    .ZN(_3984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8912_ (.A1(_3981_),
    .A2(_1100_),
    .B(_3984_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8913_ (.A1(\as2650.stack[2][6] ),
    .A2(_3982_),
    .ZN(_3985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8914_ (.A1(_3981_),
    .A2(_1108_),
    .B(_3985_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8915_ (.A1(\as2650.stack[2][7] ),
    .A2(_3982_),
    .ZN(_3986_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8916_ (.A1(_3981_),
    .A2(_1115_),
    .B(_3986_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8917_ (.A1(_2171_),
    .A2(_1687_),
    .ZN(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8918_ (.A1(_3047_),
    .A2(_1687_),
    .B(_3987_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8919_ (.A1(_2176_),
    .A2(_1686_),
    .ZN(_3988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8920_ (.A1(_1632_),
    .A2(_1687_),
    .B(_3988_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8921_ (.A1(_1513_),
    .A2(_2120_),
    .A3(_2991_),
    .A4(_1576_),
    .ZN(_3989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8922_ (.A1(_2601_),
    .A2(_1412_),
    .B(_1432_),
    .ZN(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8923_ (.A1(_1189_),
    .A2(_0696_),
    .B(_3990_),
    .ZN(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8924_ (.A1(_1435_),
    .A2(_2270_),
    .ZN(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8925_ (.A1(_1486_),
    .A2(_2198_),
    .ZN(_3993_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8926_ (.A1(_1155_),
    .A2(_3647_),
    .ZN(_3994_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _8927_ (.A1(_4202_),
    .A2(_3994_),
    .A3(_1478_),
    .A4(_1463_),
    .ZN(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8928_ (.A1(_3992_),
    .A2(_3993_),
    .A3(_2921_),
    .A4(_3995_),
    .ZN(_3996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8929_ (.A1(_1378_),
    .A2(_1477_),
    .ZN(_3997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8930_ (.A1(_1607_),
    .A2(_1420_),
    .B(_1398_),
    .ZN(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8931_ (.A1(_3997_),
    .A2(_3998_),
    .ZN(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _8932_ (.A1(_4234_),
    .A2(_1455_),
    .A3(_1370_),
    .A4(_1408_),
    .Z(_4000_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8933_ (.A1(_2136_),
    .A2(_1403_),
    .A3(_1371_),
    .ZN(_4001_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8934_ (.A1(_4312_),
    .A2(_2207_),
    .B1(_4000_),
    .B2(_2194_),
    .C(_4001_),
    .ZN(_4002_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _8935_ (.A1(_1564_),
    .A2(_2235_),
    .A3(_2254_),
    .A4(_4002_),
    .Z(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _8936_ (.A1(_3991_),
    .A2(_3996_),
    .A3(_3999_),
    .A4(_4003_),
    .ZN(_4004_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8937_ (.A1(_3989_),
    .A2(_4004_),
    .Z(_4005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8938_ (.I(_1503_),
    .ZN(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8939_ (.A1(_0624_),
    .A2(_4006_),
    .B(_1499_),
    .ZN(_4007_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8940_ (.A1(_0879_),
    .A2(_0875_),
    .B(_0872_),
    .C(_0536_),
    .ZN(_4008_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8941_ (.A1(_0620_),
    .A2(_4007_),
    .B(_4008_),
    .ZN(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8942_ (.A1(_2588_),
    .A2(_4298_),
    .A3(_4009_),
    .ZN(_4010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8943_ (.A1(_3719_),
    .A2(_3001_),
    .ZN(_4011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8944_ (.A1(_4354_),
    .A2(_3010_),
    .B(_1578_),
    .ZN(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8945_ (.A1(_3719_),
    .A2(_1636_),
    .B1(_4011_),
    .B2(_4012_),
    .C(_1575_),
    .ZN(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8946_ (.A1(_3718_),
    .A2(_4398_),
    .B(_4013_),
    .C(_2317_),
    .ZN(_4014_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8947_ (.A1(_4010_),
    .A2(_4014_),
    .A3(_4005_),
    .ZN(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8948_ (.A1(\as2650.carry ),
    .A2(_4005_),
    .B(_4015_),
    .ZN(_4016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8949_ (.A1(_3638_),
    .A2(_4016_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8950_ (.A1(_2999_),
    .A2(_1412_),
    .ZN(_4017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8951_ (.A1(_1683_),
    .A2(_4017_),
    .ZN(_4018_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8952_ (.A1(_4494_),
    .A2(_3331_),
    .Z(_4019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8953_ (.A1(_0439_),
    .A2(_0972_),
    .ZN(_4020_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8954_ (.A1(_0972_),
    .A2(_4019_),
    .B(_4020_),
    .C(_4466_),
    .ZN(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8955_ (.A1(_4466_),
    .A2(_4499_),
    .B(_4021_),
    .C(_2226_),
    .ZN(_4022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8956_ (.A1(_4018_),
    .A2(_4022_),
    .ZN(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8957_ (.A1(_4490_),
    .A2(_3444_),
    .B1(_4019_),
    .B2(_3047_),
    .ZN(_4024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8958_ (.A1(_3078_),
    .A2(_4023_),
    .B(_4024_),
    .ZN(_4025_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8959_ (.A1(_2999_),
    .A2(_1363_),
    .A3(_1399_),
    .A4(_1405_),
    .ZN(_4026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8960_ (.A1(_1365_),
    .A2(_1390_),
    .ZN(_4027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _8961_ (.A1(_4026_),
    .A2(_4027_),
    .B(_2222_),
    .ZN(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8962_ (.A1(_1624_),
    .A2(_1381_),
    .A3(_1357_),
    .ZN(_4029_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _8963_ (.A1(_4393_),
    .A2(_2253_),
    .A3(_3992_),
    .A4(_1474_),
    .Z(_4030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8964_ (.A1(_1188_),
    .A2(_2292_),
    .B(_2242_),
    .ZN(_4031_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _8965_ (.A1(_3724_),
    .A2(_2344_),
    .A3(_1383_),
    .A4(_4031_),
    .ZN(_4032_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8966_ (.A1(_2274_),
    .A2(_4029_),
    .A3(_4030_),
    .A4(_4032_),
    .ZN(_4033_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8967_ (.A1(_0408_),
    .A2(_3182_),
    .A3(_2142_),
    .A4(_2694_),
    .ZN(_4034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8968_ (.A1(_3068_),
    .A2(_0952_),
    .ZN(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8969_ (.A1(_2221_),
    .A2(_3182_),
    .A3(_0941_),
    .ZN(_4036_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8970_ (.A1(_1433_),
    .A2(_4034_),
    .A3(_4035_),
    .A4(_4036_),
    .ZN(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8971_ (.A1(_1351_),
    .A2(_1374_),
    .A3(_2193_),
    .ZN(_4038_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8972_ (.A1(_2949_),
    .A2(_3152_),
    .A3(_4038_),
    .ZN(_4039_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _8973_ (.A1(_4028_),
    .A2(_4033_),
    .A3(_4037_),
    .A4(_4039_),
    .ZN(_4040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8974_ (.A1(_1683_),
    .A2(_2195_),
    .B(_4040_),
    .ZN(_4041_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8975_ (.I0(_4025_),
    .I1(_1048_),
    .S(_4041_),
    .Z(_4042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8976_ (.A1(_3638_),
    .A2(_4042_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8977_ (.A1(_1680_),
    .A2(_2195_),
    .B(_4040_),
    .ZN(_4043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8978_ (.A1(_1551_),
    .A2(_4017_),
    .ZN(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8979_ (.A1(_0330_),
    .A2(_0971_),
    .ZN(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8980_ (.A1(_0382_),
    .A2(_0971_),
    .B(_4045_),
    .C(_1187_),
    .ZN(_4046_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8981_ (.A1(_4466_),
    .A2(_0491_),
    .B(_4046_),
    .C(_1624_),
    .ZN(_4047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8982_ (.A1(_4044_),
    .A2(_4047_),
    .B(_2192_),
    .ZN(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8983_ (.A1(_0492_),
    .A2(_2192_),
    .B(_4048_),
    .C(_3062_),
    .ZN(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8984_ (.A1(_3114_),
    .A2(_0492_),
    .B(_4049_),
    .ZN(_4050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8985_ (.A1(_4043_),
    .A2(_4050_),
    .ZN(_4051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8986_ (.A1(_1046_),
    .A2(_4043_),
    .B(_4051_),
    .ZN(_4052_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8987_ (.A1(_2231_),
    .A2(_4052_),
    .Z(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8988_ (.I(_4053_),
    .Z(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8989_ (.A1(_1669_),
    .A2(_2195_),
    .B(_4040_),
    .ZN(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8990_ (.A1(_1478_),
    .A2(_3503_),
    .Z(_4055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8991_ (.A1(_1669_),
    .A2(_4017_),
    .ZN(_4056_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8992_ (.A1(_4503_),
    .A2(_3009_),
    .A3(_4467_),
    .A4(_0972_),
    .ZN(_4057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8993_ (.A1(_4056_),
    .A2(_4057_),
    .B(_3503_),
    .ZN(_4058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8994_ (.A1(_0495_),
    .A2(_4055_),
    .B(_4058_),
    .C(_4054_),
    .ZN(_4059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8995_ (.A1(_0495_),
    .A2(_4054_),
    .B(_4059_),
    .C(_3970_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _8996_ (.A1(_1411_),
    .A2(_1398_),
    .A3(_1524_),
    .B(_4004_),
    .ZN(_4060_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8997_ (.A1(_1578_),
    .A2(_1421_),
    .B(_3022_),
    .C(_1520_),
    .ZN(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8998_ (.A1(_3762_),
    .A2(_4061_),
    .ZN(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8999_ (.A1(_3718_),
    .A2(_4062_),
    .ZN(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9000_ (.A1(_3718_),
    .A2(_1539_),
    .B(_4063_),
    .ZN(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _9001_ (.A1(_4334_),
    .A2(_0621_),
    .Z(_4065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9002_ (.A1(_0633_),
    .A2(_4065_),
    .B(_2587_),
    .ZN(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9003_ (.A1(_0634_),
    .A2(_4065_),
    .B(_4066_),
    .ZN(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _9004_ (.A1(_2215_),
    .A2(_4064_),
    .B(_4060_),
    .C(_4067_),
    .ZN(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _9005_ (.A1(_1602_),
    .A2(_4060_),
    .B(_4068_),
    .C(_3970_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _9006_ (.A1(_1553_),
    .A2(_1524_),
    .B(_1433_),
    .C(_3997_),
    .ZN(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _9007_ (.A1(_3991_),
    .A2(_3996_),
    .A3(_4003_),
    .A4(_4069_),
    .ZN(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _9008_ (.I0(_0871_),
    .I1(_0872_),
    .S(_0883_),
    .Z(_4071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9009_ (.A1(_1383_),
    .A2(_3011_),
    .ZN(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _9010_ (.A1(_2317_),
    .A2(_3012_),
    .A3(_4072_),
    .ZN(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _9011_ (.A1(_2215_),
    .A2(_4071_),
    .B(_4073_),
    .C(_4070_),
    .ZN(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9012_ (.A1(\as2650.overflow ),
    .A2(_4070_),
    .B(_4074_),
    .ZN(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9013_ (.A1(_3638_),
    .A2(_4075_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9014_ (.A1(_1404_),
    .A2(_2300_),
    .ZN(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _9015_ (.A1(_1695_),
    .A2(_1522_),
    .B(_0655_),
    .C(_2288_),
    .ZN(_4077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9016_ (.A1(_2993_),
    .A2(_1371_),
    .B(_2412_),
    .ZN(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9017_ (.A1(_4077_),
    .A2(_4078_),
    .ZN(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _9018_ (.A1(_3043_),
    .A2(_4076_),
    .B(_4079_),
    .ZN(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9019_ (.A1(_3018_),
    .A2(_4080_),
    .ZN(_4081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9020_ (.A1(_3058_),
    .A2(_1383_),
    .ZN(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9021_ (.A1(_3019_),
    .A2(_4082_),
    .ZN(_4083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9022_ (.A1(_4442_),
    .A2(_4081_),
    .ZN(_4084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _9023_ (.A1(_4081_),
    .A2(_4083_),
    .B(_4084_),
    .C(_3118_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9024_ (.A1(_3015_),
    .A2(_4080_),
    .ZN(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9025_ (.A1(_3016_),
    .A2(_4082_),
    .ZN(_4086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9026_ (.A1(_4357_),
    .A2(_4085_),
    .ZN(_4087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _9027_ (.A1(_4085_),
    .A2(_4086_),
    .B(_4087_),
    .C(_3118_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9028_ (.A1(_3005_),
    .A2(_4080_),
    .B(_1492_),
    .ZN(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _9029_ (.I(_4080_),
    .ZN(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _9030_ (.A1(_3006_),
    .A2(_4089_),
    .A3(_4082_),
    .ZN(_4090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9031_ (.A1(_4088_),
    .A2(_4090_),
    .B(_1428_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9032_ (.A1(_0793_),
    .A2(_1417_),
    .ZN(_4091_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _9033_ (.A1(_1689_),
    .A2(_3058_),
    .A3(_1413_),
    .ZN(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _9034_ (.A1(_3009_),
    .A2(_4515_),
    .A3(_1405_),
    .A4(_2300_),
    .ZN(_4093_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _9035_ (.A1(_2199_),
    .A2(_1695_),
    .A3(_1468_),
    .A4(_4167_),
    .Z(_4094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9036_ (.A1(_4078_),
    .A2(_4094_),
    .ZN(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9037_ (.A1(_4093_),
    .A2(_4095_),
    .ZN(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9038_ (.A1(_4091_),
    .A2(_4092_),
    .B(_4096_),
    .ZN(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9039_ (.A1(_3024_),
    .A2(_4096_),
    .B(_1583_),
    .ZN(_4098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9040_ (.A1(_2231_),
    .A2(_4098_),
    .ZN(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9041_ (.A1(_4097_),
    .A2(_4099_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9042_ (.A1(_3018_),
    .A2(_4096_),
    .B(\as2650.psu[4] ),
    .ZN(_4100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9043_ (.A1(_4515_),
    .A2(_1402_),
    .ZN(_4101_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _9044_ (.A1(_3097_),
    .A2(_4101_),
    .A3(_4076_),
    .B(_4095_),
    .ZN(_4102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9045_ (.A1(_3058_),
    .A2(_1413_),
    .B(_4102_),
    .ZN(_4103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9046_ (.A1(_3019_),
    .A2(_4103_),
    .ZN(_4104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9047_ (.A1(_4100_),
    .A2(_4104_),
    .B(_1428_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9048_ (.A1(_3015_),
    .A2(_4096_),
    .B(\as2650.psu[3] ),
    .ZN(_4105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9049_ (.A1(_3016_),
    .A2(_4103_),
    .ZN(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9050_ (.A1(_4105_),
    .A2(_4106_),
    .B(_1428_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9051_ (.D(_0000_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9052_ (.D(_0001_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9053_ (.D(_0002_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9054_ (.D(_0003_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9055_ (.D(_0004_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9056_ (.D(_0005_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.r123[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9057_ (.D(_0006_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9058_ (.D(_0007_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9059_ (.D(_0008_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9060_ (.D(_0009_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9061_ (.D(_0010_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9062_ (.D(_0011_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9063_ (.D(_0012_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9064_ (.D(_0013_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9065_ (.D(_0014_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9066_ (.D(_0015_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9067_ (.D(_0016_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9068_ (.D(_0017_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9069_ (.D(_0018_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9070_ (.D(_0019_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9071_ (.D(_0020_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9072_ (.D(_0021_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9073_ (.D(_0022_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9074_ (.D(_0023_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9075_ (.D(_0024_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9076_ (.D(_0025_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9077_ (.D(_0026_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9078_ (.D(_0027_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9079_ (.D(_0028_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9080_ (.D(_0029_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9081_ (.D(_0030_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9082_ (.D(_0031_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.r123_2[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9083_ (.D(_0032_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.r123_2[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9084_ (.D(_0033_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.r123_2[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9085_ (.D(_0034_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.r123_2[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9086_ (.D(_0035_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.r123_2[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9087_ (.D(_0036_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.r123_2[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9088_ (.D(_0037_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.r123_2[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9089_ (.D(_0038_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.r123_2[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9090_ (.D(_0039_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9091_ (.D(_0040_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9092_ (.D(_0041_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9093_ (.D(_0042_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9094_ (.D(_0043_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9095_ (.D(_0044_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9096_ (.D(_0045_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9097_ (.D(_0046_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9098_ (.D(_0047_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9099_ (.D(_0048_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9100_ (.D(_0049_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9101_ (.D(_0050_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9102_ (.D(_0051_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9103_ (.D(_0052_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9104_ (.D(_0053_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9105_ (.D(_0054_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9106_ (.D(_0055_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9107_ (.D(_0056_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9108_ (.D(_0057_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9109_ (.D(_0058_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9110_ (.D(_0059_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9111_ (.D(_0060_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9112_ (.D(_0061_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9113_ (.D(_0062_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9114_ (.D(_0063_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9115_ (.D(_0064_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9116_ (.D(_0065_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9117_ (.D(_0066_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9118_ (.D(_0067_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.alu_op[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9119_ (.D(_0068_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.alu_op[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9120_ (.D(_0069_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\as2650.alu_op[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9121_ (.D(_0070_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123_2[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9122_ (.D(_0071_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123_2[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9123_ (.D(_0072_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123_2[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9124_ (.D(_0073_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.r123_2[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9125_ (.D(_0074_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.r123_2[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9126_ (.D(_0075_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.r123_2[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9127_ (.D(_0076_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.r123_2[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9128_ (.D(_0077_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123_2[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9129_ (.D(_0078_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9130_ (.D(_0079_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9131_ (.D(_0080_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9132_ (.D(_0081_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9133_ (.D(_0082_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9134_ (.D(_0083_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9135_ (.D(_0084_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9136_ (.D(_0085_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9137_ (.D(_0086_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9138_ (.D(_0087_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9139_ (.D(_0088_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9140_ (.D(_0089_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9141_ (.D(_0090_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9142_ (.D(_0091_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9143_ (.D(_0092_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9144_ (.D(_0093_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.r123[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9145_ (.D(_0094_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.r123[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9146_ (.D(_0095_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.r123[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9147_ (.D(_0096_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.r123[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9148_ (.D(_0097_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.r123[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9149_ (.D(_0098_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.r123[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9150_ (.D(_0099_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.r123[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9151_ (.D(_0100_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.r123[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9152_ (.D(_0101_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9153_ (.D(_0102_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9154_ (.D(_0103_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9155_ (.D(_0104_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9156_ (.D(_0105_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9157_ (.D(_0106_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9158_ (.D(_0107_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9159_ (.D(_0108_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9160_ (.D(_0109_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123_2[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9161_ (.D(_0110_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123_2[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9162_ (.D(_0111_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123_2[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9163_ (.D(_0112_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123_2[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9164_ (.D(_0113_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123_2[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9165_ (.D(_0114_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123_2[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9166_ (.D(_0115_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123_2[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9167_ (.D(_0116_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.r123_2[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9168_ (.D(_0117_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9169_ (.D(_0118_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9170_ (.D(_0119_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9171_ (.D(_0120_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9172_ (.D(_0121_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9173_ (.D(_0122_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9174_ (.D(_0123_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9175_ (.D(_0124_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9176_ (.D(_0125_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9177_ (.D(_0126_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9178_ (.D(_0127_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9179_ (.D(_0128_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9180_ (.D(_0129_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9181_ (.D(_0130_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.addr_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9182_ (.D(_0131_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.addr_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9183_ (.D(_0132_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9184_ (.D(_0133_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9185_ (.D(_0134_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9186_ (.D(_0135_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9187_ (.D(_0136_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9188_ (.D(_0137_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9189_ (.D(_0138_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9190_ (.D(_0139_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9191_ (.D(_0140_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9192_ (.D(_0141_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9193_ (.D(_0142_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(net34));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9194_ (.D(_0143_),
    .CLK(clknet_opt_3_0_wb_clk_i),
    .Q(net35));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9195_ (.D(_0144_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(net36));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9196_ (.D(_0145_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(net37));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9197_ (.D(_0146_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(net38));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9198_ (.D(_0147_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(net39));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9199_ (.D(_0148_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(net40));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9200_ (.D(_0149_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9201_ (.D(_0150_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9202_ (.D(_0151_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.idx_ctrl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9203_ (.D(_0152_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.idx_ctrl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9204_ (.D(_0153_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.holding_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9205_ (.D(_0154_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9206_ (.D(_0155_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9207_ (.D(_0156_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9208_ (.D(_0157_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9209_ (.D(_0158_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9210_ (.D(_0159_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9211_ (.D(_0160_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9212_ (.D(_0161_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9213_ (.D(_0162_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9214_ (.D(_0163_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9215_ (.D(_0164_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9216_ (.D(_0165_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _9217_ (.D(_0166_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9218_ (.D(_0167_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\as2650.cycle[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9219_ (.D(_0168_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9220_ (.D(_0169_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9221_ (.D(_0170_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9222_ (.D(_0171_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9223_ (.D(_0172_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9224_ (.D(_0173_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9225_ (.D(_0174_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9226_ (.D(_0175_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9227_ (.D(_0176_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9228_ (.D(_0177_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9229_ (.D(_0178_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9230_ (.D(_0179_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9231_ (.D(_0180_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9232_ (.D(_0181_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9233_ (.D(_0182_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9234_ (.D(_0183_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9235_ (.D(_0184_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.pc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9236_ (.D(_0185_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.pc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9237_ (.D(_0186_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9238_ (.D(_0187_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9239_ (.D(_0188_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9240_ (.D(_0189_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9241_ (.D(_0190_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9242_ (.D(_0191_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9243_ (.D(_0192_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9244_ (.D(_0193_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9245_ (.D(_0194_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9246_ (.D(_0195_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9247_ (.D(_0196_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9248_ (.D(_0197_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9249_ (.D(_0198_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9250_ (.D(_0199_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9251_ (.D(_0200_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9252_ (.D(_0201_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9253_ (.D(_0202_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9254_ (.D(_0203_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9255_ (.D(_0204_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9256_ (.D(_0205_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9257_ (.D(_0206_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9258_ (.D(_0207_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9259_ (.D(_0208_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9260_ (.D(_0209_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9261_ (.D(_0210_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9262_ (.D(_0211_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9263_ (.D(_0212_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9264_ (.D(_0213_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9265_ (.D(_0214_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9266_ (.D(_0215_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9267_ (.D(_0216_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9268_ (.D(_0217_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9269_ (.D(_0218_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9270_ (.D(_0219_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9271_ (.D(_0220_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9272_ (.D(_0221_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9273_ (.D(_0222_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9274_ (.D(_0223_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9275_ (.D(_0224_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9276_ (.D(_0225_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9277_ (.D(_0226_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9278_ (.D(_0227_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9279_ (.D(_0228_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9280_ (.D(_0229_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9281_ (.D(_0230_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9282_ (.D(_0231_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9283_ (.D(_0232_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9284_ (.D(_0233_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9285_ (.D(_0234_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9286_ (.D(_0235_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9287_ (.D(_0236_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9288_ (.D(_0237_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9289_ (.D(_0238_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.r123[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9290_ (.D(_0239_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.r123[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9291_ (.D(_0240_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9292_ (.D(_0241_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.r123[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9293_ (.D(_0242_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.r123[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9294_ (.D(_0243_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.r123[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9295_ (.D(_0244_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.r123[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9296_ (.D(_0245_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9297_ (.D(_0246_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9298_ (.D(_0247_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9299_ (.D(_0248_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9300_ (.D(_0249_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9301_ (.D(_0250_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9302_ (.D(_0251_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.r123[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9303_ (.D(_0252_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9304_ (.D(_0253_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9305_ (.D(_0254_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(net41));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9306_ (.D(_0255_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(net42));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9307_ (.D(_0256_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(net43));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9308_ (.D(_0257_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(net44));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9309_ (.D(_0258_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(net45));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9310_ (.D(_0259_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9311_ (.D(_0260_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9312_ (.D(_0261_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9313_ (.D(_0262_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9314_ (.D(_0263_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9315_ (.D(_0264_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9316_ (.D(_0265_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9317_ (.D(_0266_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9318_ (.D(_0267_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9319_ (.D(_0268_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9320_ (.D(_0269_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9321_ (.D(_0270_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9322_ (.D(_0271_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9323_ (.D(_0272_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.carry ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9324_ (.D(_0273_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9325_ (.D(_0274_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9326_ (.D(_0275_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.psu[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9327_ (.D(_0276_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9328_ (.D(_0277_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9329_ (.D(_0278_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9330_ (.D(_0279_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9331_ (.D(_0280_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9332_ (.D(_0281_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9333_ (.D(_0282_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9334_ (.D(_0283_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_86 (.Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_87 (.Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_88 (.Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_89 (.Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_90 (.Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_91 (.Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_92 (.Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_93 (.Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_94 (.Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_95 (.Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_56 (.ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_57 (.ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_58 (.ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_59 (.ZN(net59));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_60 (.ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_61 (.ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_62 (.ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_63 (.ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_64 (.ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_65 (.ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_66 (.ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_67 (.ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_68 (.ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_69 (.ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_70 (.ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_71 (.ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_85 (.Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9376_ (.I(net46),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9377_ (.I(net46),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9378_ (.I(net46),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9379_ (.I(net48),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9380_ (.I(net46),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9381_ (.I(net47),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9382_ (.I(net48),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(io_in[10]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input2 (.I(io_in[11]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(io_in[12]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(io_in[13]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input5 (.I(io_in[33]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(io_in[5]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input7 (.I(io_in[6]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input8 (.I(io_in[7]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input9 (.I(io_in[8]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input10 (.I(io_in[9]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output11 (.I(net11),
    .Z(io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output12 (.I(net12),
    .Z(io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output13 (.I(net47),
    .Z(io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output14 (.I(net14),
    .Z(io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output15 (.I(net15),
    .Z(io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output16 (.I(net16),
    .Z(io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output17 (.I(net17),
    .Z(io_oeb[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output18 (.I(net18),
    .Z(io_oeb[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output19 (.I(net19),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output20 (.I(net20),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output21 (.I(net21),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output22 (.I(net22),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output23 (.I(net23),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output24 (.I(net24),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output25 (.I(net25),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output26 (.I(net26),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output27 (.I(net27),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output28 (.I(net28),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output29 (.I(net29),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output30 (.I(net30),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output31 (.I(net31),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output32 (.I(net32),
    .Z(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output33 (.I(net33),
    .Z(io_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output34 (.I(net34),
    .Z(io_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output35 (.I(net35),
    .Z(io_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output36 (.I(net36),
    .Z(io_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output37 (.I(net37),
    .Z(io_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output38 (.I(net38),
    .Z(io_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output39 (.I(net39),
    .Z(io_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output40 (.I(net40),
    .Z(io_out[32]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output41 (.I(net41),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output42 (.I(net42),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output43 (.I(net43),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output44 (.I(net44),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output45 (.I(net45),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout46 (.I(net48),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout47 (.I(net48),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout48 (.I(net13),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout49 (.I(net25),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout50 (.I(net26),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout51 (.I(net40),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout52 (.I(net38),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout53 (.I(net31),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout54 (.I(net28),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_55 (.ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.I(clknet_3_2__leaf_wb_clk_i),
    .Z(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.I(clknet_3_2__leaf_wb_clk_i),
    .Z(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.I(clknet_3_3__leaf_wb_clk_i),
    .Z(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_8_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_10_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.I(clknet_3_3__leaf_wb_clk_i),
    .Z(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.I(clknet_3_2__leaf_wb_clk_i),
    .Z(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.I(clknet_3_2__leaf_wb_clk_i),
    .Z(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.I(clknet_3_2__leaf_wb_clk_i),
    .Z(clknet_leaf_16_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.I(clknet_3_2__leaf_wb_clk_i),
    .Z(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.I(clknet_opt_2_0_wb_clk_i),
    .Z(clknet_leaf_19_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_22_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_wb_clk_i (.I(clknet_opt_5_0_wb_clk_i),
    .Z(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_wb_clk_i (.I(clknet_opt_4_0_wb_clk_i),
    .Z(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_wb_clk_i (.I(clknet_opt_1_0_wb_clk_i),
    .Z(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_0__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_1__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_2__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_3__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_4__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_5__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_6__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_7__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_1_0_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_opt_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_2_0_wb_clk_i (.I(clknet_3_3__leaf_wb_clk_i),
    .Z(clknet_opt_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_3_0_wb_clk_i (.I(clknet_3_3__leaf_wb_clk_i),
    .Z(clknet_opt_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_4_0_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_opt_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_5_0_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_opt_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9107__D (.I(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9118__D (.I(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9119__D (.I(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9120__D (.I(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9186__D (.I(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9203__D (.I(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9216__D (.I(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9227__D (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9229__D (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9230__D (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9238__D (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9239__D (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9240__D (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9241__D (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9243__D (.I(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9329__D (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__A1 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__A1 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__A1 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__I (.I(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__A2 (.I(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A2 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__A1 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__I (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__A2 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__A2 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__A2 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A1 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__A1 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__A1 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__I (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__A1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__A1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__C (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__A2 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__A2 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__A2 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A1 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__A2 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__A2 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__A2 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__A2 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__B (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A2 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__A1 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__C (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__A2 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__C (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__S (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__C (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__C (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__C (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8534__A2 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__A1 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5954__A1 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__A2 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__A1 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__A1 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__A1 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__A1 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__A2 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__I (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__A2 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__A2 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__C (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__A2 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__B (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8533__A2 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7188__A2 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__A1 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__A2 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__B2 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__B2 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__B2 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__A2 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__C (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__B (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8532__A2 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7194__A2 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5951__A1 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__A2 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__B2 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6483__A1 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__A1 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__I (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8979__A1 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6244__A2 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__A1 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__I (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6439__A1 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__I (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__A1 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__A1 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8506__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__I (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__I (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7922__A3 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7057__A2 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6993__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__A2 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8782__A3 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__B2 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__A3 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__A3 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__S1 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__S (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__S1 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__S (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8153__A2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8108__A2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__A2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__B1 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__A1 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__A2 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__A1 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__I (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__B2 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__B2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__A2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__A3 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__A2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__A3 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__A1 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__A2 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5008__I (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__A1 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__I (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8537__I (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__A2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__A2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8109__A1 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7278__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7258__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__I (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7240__A1 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6322__A2 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__I (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__I (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8053__A1 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7194__A1 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__B2 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__I (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8060__A1 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8054__A1 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7188__A1 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__I (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7212__B2 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6405__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__A1 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__A1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__A3 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__B2 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__A2 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__A1 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__A1 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__I (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__A3 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8546__A1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7090__A2 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__B2 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__A2 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8542__A2 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__A2 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__B2 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__I (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8857__A1 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8525__A1 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5948__A1 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8828__A1 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8796__A1 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__A2 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8210__B2 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8165__I (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8074__B2 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__A1 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8245__B1 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8075__I (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8033__I (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__A2 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8276__A1 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__I (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__I (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__I (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8980__A1 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__A1 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__A1 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__A1 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8306__B2 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8168__A1 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8028__A1 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__I (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__A1 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__I (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__A1 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__A1 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8243__B2 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8162__I (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8078__B2 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__I (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8306__A1 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8028__B2 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__I (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__I (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5512__A2 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__A1 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__A2 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__A2 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__I (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__B2 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__B2 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__B2 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8366__A1 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__A1 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__A2 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__B (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7900__A1 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__A1 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__A3 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__A1 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7078__I (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6914__A1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__A1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8232__A2 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8184__A2 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8113__I (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5070__I (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8967__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8000__A2 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7211__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__I (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7938__A2 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7923__A1 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7567__A1 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__A4 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__A1 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__A1 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__B (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5189__A1 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__B1 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__A1 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__A1 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__A1 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__A1 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__I (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__A1 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__I (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__A2 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__A2 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__A2 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__I (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__A2 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__A2 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__I (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__A2 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__A1 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__A1 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__B1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__B (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__A2 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__A2 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__A2 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__B (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__B2 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__B2 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__A1 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__C (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__B (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__A1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__B2 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__A1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__B2 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8552__A2 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__A2 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__A1 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__A2 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__A1 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6244__A1 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__I (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__I (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8953__A1 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7826__A1 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__I (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__A1 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8862__A1 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8501__A2 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__B1 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__A2 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6777__A1 (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6751__A1 (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6534__A1 (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__I (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6750__B2 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__A1 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__I (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__A1 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8188__A2 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8187__A2 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8155__A2 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__A2 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__A2 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5112__A2 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__A2 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__A4 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__A2 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__I (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__B1 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__A2 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__A2 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__I (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__A1 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__A1 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__I (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__A2 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8153__A1 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8108__A1 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7314__A2 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__I (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7304__A1 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7249__A1 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6325__I (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5117__I (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7242__A1 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__A1 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6307__C2 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__I (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__A1 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6267__I (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__A1 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__A1 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__A2 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__A1 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__A1 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__I (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5947__A1 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__A1 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__A2 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__A1 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__B (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8564__B2 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7090__A3 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__A1 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5126__A2 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__A2 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__A2 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7304__A2 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7249__A2 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__I (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8551__A2 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__A2 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__I0 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__A2 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__A1 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__I (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__A1 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__A1 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5434__A1 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__B2 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__B2 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8550__A2 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7242__A2 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__A1 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__A2 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8831__A1 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8800__A1 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A2 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8981__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__A1 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__A1 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__I (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8984__A2 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8983__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8122__A1 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8071__A1 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8037__A1 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__I (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8277__A1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8163__A1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__I (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__I (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8995__A1 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8994__A1 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__A1 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A1 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__A1 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__B2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__B2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__B2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8308__C (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8124__B (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8039__B (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__I (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__C (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__C (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__C (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__C (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8390__A1 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5959__A1 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8867__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__B (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5675__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__A1 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__I (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__A2 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7834__A1 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__A1 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__A2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__A3 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__I (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5300__A2 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__A2 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__I (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__A2 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__A2 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__A2 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__A2 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6223__A4 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__B (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__B1 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__A1 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8940__C (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__A1 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__A1 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__B2 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8583__A2 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6204__A2 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5992__A1 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__A2 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7830__I (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__A1 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__I (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__A1 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6778__A1 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__A1 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__I (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__A1 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8222__A2 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8221__A2 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8186__A2 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__A2 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__A2 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__A2 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__A2 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__A2 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__B (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__A2 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__I (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8878__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__A2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5984__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__A2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8188__A1 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8187__A1 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7343__I (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__I (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7359__A2 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__A2 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6269__I (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__I (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__A1 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7301__A1 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__A1 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__A1 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8595__A2 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__A2 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__B (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__A1 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__A1 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5300__A1 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__A1 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__B1 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8580__B2 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7090__A4 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5982__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__A2 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__A2 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__A1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__A1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A2 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__A2 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A2 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__A1 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__B1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__A2 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__B1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__A2 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__B1 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__A2 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7351__A2 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7350__A2 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__I (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8582__A2 (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__A2 (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__A1 (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__A2 (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__B2 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__B2 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__B2 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__A1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__C (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8581__A2 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__A2 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8834__A1 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8804__A1 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__A2 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A1 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__A1 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__A1 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__A1 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__A1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__A1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__A1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__B2 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5443__B2 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__B2 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__B2 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__A2 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__A2 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__A2 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__A2 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5443__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8415__A1 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__A1 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__A2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8872__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5977__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__B (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5453__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__A4 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__I (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__A3 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__I (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__A2 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6809__A1 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__A1 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__A1 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__I (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__A1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__A1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__I (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__A1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__A2 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__A2 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__I (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8941__A1 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__B2 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__A1 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__A1 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9001__A2 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__A1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__A2 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__A1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8939__A1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5290__A2 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__A2 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__A1 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__A2 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9002__A1 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6204__A3 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5298__I (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9003__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8588__A2 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6007__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__A2 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8613__A2 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__I (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A1 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A1 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__A2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__A2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__A2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5304__I (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6255__A2 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__A4 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__B1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__B1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7433__A2 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7432__A2 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__I (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8587__A2 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__A2 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__A1 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__A2 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6768__A1 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__A3 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__I (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__A1 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__A2 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__I (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6830__A2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__B1 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__I (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__A2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6708__A1 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6580__A1 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__I (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__I (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8620__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5432__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8266__A2 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8265__A2 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8224__A2 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__A2 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9015__B (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7068__A3 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__A3 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__A1 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5675__A1 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5674__A1 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5412__S (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__A1 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__A2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__A2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__I (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__A3 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__A3 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__A2 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__I (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__S (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__A2 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__A2 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__I (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7089__A1 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__A2 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__A1 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__I (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__B1 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__A1 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6000__A1 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__I (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8597__I (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6255__A3 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__A2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__A2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5566__A1 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__A1 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__A1 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A1 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5424__A2 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__A1 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__B1 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__A2 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5424__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__B2 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8589__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7091__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5999__B2 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__A2 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8222__A1 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8221__A1 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7358__A2 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__I (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7411__A2 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__B1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__I (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__I (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8186__A1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__A1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6307__B1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__I (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8196__A1 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6965__I (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6273__I (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__A1 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8871__A1 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8580__A1 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8562__A2 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__A2 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7426__A2 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7425__A2 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__I (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8586__A2 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7353__A2 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__A1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__A2 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8839__A1 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8809__A1 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__A2 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__A1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__I (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__A1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6407__A1 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__A1 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A2 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__A2 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6090__I (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__A1 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8923__A2 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__A3 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__A2 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__A2 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__A1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__A2 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8788__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__C (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8879__A1 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__A1 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__I (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__A1 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__A1 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__B (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8437__A1 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__A2 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__A1 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__A3 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__B (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6810__A1 (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6784__A1 (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__A1 (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5381__I (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6835__A1 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__A1 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5447__I (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__A1 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__A2 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__A2 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5393__A1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__A2 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__B (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__A2 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__A1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8607__A2 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__A1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6022__A1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__I0 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7423__A2 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__I (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8604__A2 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7453__A2 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__A1 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__A2 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8601__A1 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8577__A2 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__A1 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5431__A2 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__I1 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__A1 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__A1 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__I (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8298__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8297__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8268__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5413__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__A2 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5416__A2 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5415__A2 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__A4 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5456__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__I (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5564__A2 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5563__B (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__A2 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5418__I (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__C1 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__A1 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A2 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__I (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__I (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__A1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7468__A2 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7419__A2 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6300__I (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5421__I (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7435__A1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__B1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__B2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__I (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8224__A1 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__I (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__A1 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__A1 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6014__A1 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__A2 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7460__A2 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7459__A2 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__I (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8605__A2 (.I(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7435__A2 (.I(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A1 (.I(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5437__A2 (.I(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8841__A1 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8812__A1 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5452__A2 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8442__I (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__A2 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__A2 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6860__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6730__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5448__I (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7839__A1 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__A2 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__A1 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__I (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8884__A1 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__A1 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__A1 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__A1 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5452__B (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__A2 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5484__A2 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__A2 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5458__I (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8608__A2 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6233__A2 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__A2 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9032__A1 (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6812__A1 (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__A1 (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5460__A1 (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__A3 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__A2 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__A2 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__A2 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5464__A2 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5541__A1 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__A2 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__A1 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__A1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__A2 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__A2 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__A1 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__A2 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__B (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5470__A1 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8623__A2 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__A3 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A2 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__A1 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__A2 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__A1 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7458__A2 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__I (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8622__A2 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7517__A2 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__A2 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__B2 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__I (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6030__A1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__I (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__A1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5504__A1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5491__I (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__A1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__A1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5534__A2 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__I (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__C1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__A2 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__I (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6352__I (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6255__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__A2 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8632__A1 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__A2 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__B2 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__A2 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7635__A2 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7557__A2 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7451__I (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__I (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7699__A2 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7696__A2 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7517__A1 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__I (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7595__A2 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__B1 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6240__I (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5499__I (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8268__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__A2 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5500__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7452__A2 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__I (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8621__A2 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7512__A2 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__A1 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__A2 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8844__A1 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8815__A1 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__A2 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A2 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8478__A1 (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__A1 (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__A2 (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__B (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6861__I0 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6246__B (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5576__I (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__I (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7977__A1 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__A1 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__A1 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__I (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8893__A1 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8635__A1 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__A1 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5530__A1 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__A1 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__A2 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__B1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6214__A1 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__I0 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__A1 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__A1 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9008__S (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__A2 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__A1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__I (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8817__A2 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8636__A2 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__A2 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__A2 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__B1 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__B1 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__A2 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__A2 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A2 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__A2 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__A2 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7540__A2 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__I (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8638__A2 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7519__A2 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__A2 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7532__A2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7514__A2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__I (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8637__A2 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7535__A2 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__A1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__A2 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8650__A1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__A3 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__B2 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5566__A2 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8331__A1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8330__A1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7540__A1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__I (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8300__A1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8002__I (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__I (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5569__I (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8194__A1 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8148__A2 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__I (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5570__A1 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__A1 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5572__I (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8646__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__B1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6873__B2 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6872__A1 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6054__A1 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__A1 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5582__A2 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__B2 (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8311__A1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8279__A1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8032__A1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5587__I (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8166__A1 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__A2 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__I (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A2 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__A1 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__A1 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5598__I (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__I (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__A1 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__A1 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__A1 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__A1 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7983__C (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7088__A2 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__A2 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8513__A1 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7770__I (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__A2 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__A2 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__I (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__A2 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__A1 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7866__A1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7806__I (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__A1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7011__A3 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6927__I (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6917__A1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__A2 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7778__A2 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7060__I (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__A2 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7214__A1 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__A1 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6072__B (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__A1 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__I (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__I (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__A2 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__A2 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8195__I (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7217__I (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__B1 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7519__A1 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__A2 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__I (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__B2 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7271__A2 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A1 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__A1 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A2 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7713__A2 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__A2 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7325__I (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__B (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8005__A2 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7110__A1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__I (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__A1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7123__I (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7083__A3 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__A2 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8021__I (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7758__B2 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7497__A2 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__B (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8969__A3 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__C (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__A1 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7930__A3 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6931__A1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__A1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__A1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__B (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5637__I (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__I (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__A2 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5894__I (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6116__A1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__A2 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5639__I (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__A2 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A2 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__A2 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8013__I (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7782__A1 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__I (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__A1 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7273__I (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A2 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A2 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__A2 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__A2 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__A2 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__I (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5626__I (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__A1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5673__A1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__A1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__A1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__A2 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5628__I (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__A2 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__A2 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__A2 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__I (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8497__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6439__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__A1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7980__A1 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7927__B (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__A1 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A1 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8356__A1 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8349__A1 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7595__A1 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__I (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8346__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7579__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7577__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8521__A3 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__A1 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6239__A2 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__I (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7216__A1 (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6923__A1 (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__I (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A2 (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8992__A4 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8954__A1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8953__A2 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A3 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5795__A2 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__A2 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5699__A2 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__A2 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8673__I (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__I (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6619__A1 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__A1 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__A1 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__A2 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A1 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__A1 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5695__A1 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__A2 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6579__A2 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__A2 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__I (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__A2 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__A2 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__A2 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__I (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__A3 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__A3 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__A3 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__I (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__A2 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__A3 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__A2 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__I (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8538__A2 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__A2 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__A2 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__A1 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8374__A1 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7593__A1 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__I (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8360__A1 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8357__A1 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8350__A1 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__A1 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8681__I (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__I (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6622__A1 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__A1 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A1 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__A2 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__A2 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__A2 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__A2 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5661__A2 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__A2 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5664__I (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6742__A2 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__A4 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__A4 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__I (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8558__A2 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__A4 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__A4 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5670__A1 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8395__A1 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7635__A1 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__I (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8394__A1 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8372__A1 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7649__A1 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__A1 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8685__I (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5671__I (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6624__A1 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__A1 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5850__A1 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5673__A2 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__A2 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__A2 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6483__A2 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5676__I (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__A2 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__A2 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__A2 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5677__I (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6786__A2 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__A2 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__A2 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5678__I (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8575__A2 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6801__A2 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6730__A2 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__A1 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7682__A1 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7672__A1 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__A1 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__S (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__A2 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5691__A2 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__A2 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8688__I (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__I (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6626__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__A2 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6576__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6542__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__I (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__I (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6519__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6514__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__I (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8594__A2 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__A2 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__A2 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5692__A1 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8450__A1 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8441__A1 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8423__A1 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5691__A1 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8691__I (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__I (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6628__A1 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__A1 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A1 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5695__A2 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8612__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6768__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A1 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8468__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8460__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8451__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5699__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6630__A1 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__A1 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__A1 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__A2 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8482__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8469__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8466__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7972__B2 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7900__B2 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__A1 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__A1 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8515__A1 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7059__A1 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__A3 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__A2 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__A2 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__I (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6706__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__B1 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6539__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__I (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8624__A2 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__B1 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6810__A2 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__A2 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8697__I (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__I (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A2 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8986__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6593__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8975__I1 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8896__A2 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__A2 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__A2 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8719__A2 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__A2 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__I (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__I (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__I (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5738__I (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__I (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8858__A1 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8527__B2 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__I0 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__A1 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8007__A1 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7221__A1 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7204__A1 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__I (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8011__A1 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8005__A1 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8003__A1 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5733__I (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8047__A1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8046__A1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8042__A1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5735__A1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__I (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5737__I (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8900__A2 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6597__A1 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__A1 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__A2 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8863__A1 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7817__I (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__A1 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__A1 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8089__A1 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7278__A1 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7177__I (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__I (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8087__A1 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8064__A1 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7227__A1 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__A1 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6656__I (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__I (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8902__A2 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6599__A1 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__A1 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__A2 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8142__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7314__A1 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7261__A1 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5751__I (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8143__A1 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8098__A1 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7283__A1 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__I (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8137__A1 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7287__A1 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__A1 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__A1 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6659__I (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__I (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8904__A2 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6601__A1 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__A1 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__A2 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8179__A1 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8148__A1 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8140__A1 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5762__I (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8175__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7318__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__I (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__I (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8906__A2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6603__A1 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5812__A1 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__A2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8603__A1 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7836__A1 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__I0 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8217__A1 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8216__A1 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7409__A1 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__I1 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6665__I (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__I (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8910__A2 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__A1 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__A1 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5775__A2 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7467__A1 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7419__A1 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__I (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8250__A1 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8219__A1 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7417__A1 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__A1 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6670__I (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5780__I (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8912__A2 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6609__A1 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5818__A1 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__A2 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8888__A1 (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8633__A1 (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7844__A1 (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A1 (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8254__A1 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7502__A1 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7449__I (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5785__I (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8285__A1 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8252__A1 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7469__A1 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__A1 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6673__I (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5789__I (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8914__A2 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6611__A1 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__A1 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5791__A2 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8356__A2 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7557__A1 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7492__I (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5793__I (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8317__A1 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8290__A1 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8287__A1 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5795__A1 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6676__I (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__I (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8916__A2 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6613__A1 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5822__A1 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__A2 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8700__A3 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6614__A2 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6362__A3 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5801__I (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__I (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__I (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5804__I (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5803__I (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5822__A2 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__A2 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5818__A2 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__A2 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__A2 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5819__A2 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5817__A2 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5815__A2 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__I (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__I (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__A2 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5850__A2 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A2 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__A2 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A2 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__A2 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A2 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__A2 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A2 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5851__A2 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A2 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__A2 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8518__A1 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7859__A1 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6193__B (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5861__I (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8926__A1 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8102__A1 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7330__I (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__A1 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__A1 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__A3 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__A2 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__A2 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__A3 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__A2 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5888__A2 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__A2 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5910__A2 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__A2 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__A3 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__A3 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5940__I (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__I (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__B (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5918__I (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5902__I (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__A1 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__A2 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5915__I (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__I (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__A1 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__A1 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__A1 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__A2 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5970__A2 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5934__A2 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__A1 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5877__A2 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__B (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5898__I (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__A3 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__A4 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__A2 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__C (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6679__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6060__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__B (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__C (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5996__I (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__I (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7768__B (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6153__A1 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__A2 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__I (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A2 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__A1 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__B (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A1 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__I (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8980__C (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8557__A1 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8491__A1 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__A1 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8964__A1 (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7108__A2 (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6936__A1 (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__I (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8923__A1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8296__A1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7416__I (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__A2 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__I (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5930__I (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__S (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__A2 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8521__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8519__A1 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__I (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__A1 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__I (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__I (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__I (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8559__A2 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8547__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5917__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8017__A1 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7193__A1 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6905__I (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5916__A1 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__I (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__I (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7029__A1 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6984__I (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__A2 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__A1 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__B1 (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5914__I (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6683__A1 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__A1 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__B1 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8778__A1 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8590__A1 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__A1 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__A1 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6126__A1 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__A2 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__A2 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__A2 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__A2 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5952__B (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__C (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__B1 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__C (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__I (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6953__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__A2 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6725__A1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6444__A1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__B1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8520__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7082__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__A3 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__A3 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__A2 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__A2 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__A1 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__A2 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8566__A1 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5968__A1 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5968__B (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__B (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6762__A1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5974__B1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__A2 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7344__A2 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7301__A2 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__A1 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6795__A1 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__A1 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__B1 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A2 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__A2 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6028__A2 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__A2 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A2 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__A1 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8184__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7353__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5999__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__A2 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6883__B2 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6848__A1 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6496__A1 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__B2 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__B (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__B (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__B (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__A1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6529__A1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__A2 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__B (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7726__A1 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7004__A1 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__A1 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__A1 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__A1 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6560__A1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__I (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6868__A1 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__B1 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7535__A1 (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__I (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6258__I (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__A1 (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6883__A1 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6591__A1 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6060__A3 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8555__A2 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A1 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__A3 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6072__A1 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7922__A1 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7057__B (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__A1 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__A1 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8471__A1 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7988__A1 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7966__A2 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6065__I (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8971__A1 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8012__C (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7804__I (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7808__A1 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A2 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7096__A3 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7049__A3 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__A1 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__A2 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6070__A1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7093__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__A3 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8962__A3 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7989__A1 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7093__B (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6072__A2 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7053__A1 (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__I (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__A1 (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8613__A1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6232__I (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6231__A1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__A2 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6292__I (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6122__A2 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__A1 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8506__A4 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6985__I (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__A2 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8959__A2 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7004__A2 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__A2 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__A2 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7061__A3 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__B (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__A2 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8960__A1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6145__I (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__A1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6384__A2 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6081__I (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8820__A2 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6679__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__A3 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__I (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__A1 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__A1 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__A2 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6236__I (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__A3 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8932__A3 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6294__A2 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__I (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9016__A2 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8933__A3 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__A2 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__A2 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__A1 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__A2 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A2 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__I (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8233__C (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7085__A2 (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7032__B (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__C (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8971__A2 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6154__A3 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__A2 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8778__A3 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7735__A2 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__A2 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__A1 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8643__A1 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8573__I (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8541__C (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__A2 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8929__A1 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8778__A2 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7772__B (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__A1 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7061__A2 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7052__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6094__I (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8507__C (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7236__I (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__B (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__A2 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8962__A2 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6993__A2 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__A4 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A4 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__A4 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__A3 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6126__A2 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__A2 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9020__A2 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9009__A1 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8965__A3 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__A3 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7077__I (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__A2 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__A1 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__A1 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7761__A2 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__A1 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__A2 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7730__A1 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__A2 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__I (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6102__I (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7812__I (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__I (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__A2 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__A1 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7029__A2 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__A4 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__I (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__A2 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8960__A2 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7987__A1 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__A4 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8408__A1 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7818__I (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__A1 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__A1 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__A2 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__I (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8996__A2 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8930__B (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7905__A2 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__A2 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8555__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7049__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__A2 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__A2 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__A1 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6116__A2 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9043__A2 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7866__A3 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__A1 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8933__A2 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8555__A3 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__A3 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9014__A1 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7976__A2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__A2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__A2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9034__A3 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8959__A4 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__A4 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8932__A4 (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__C (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8225__A1 (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7431__A1 (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__A2 (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__I (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8996__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6132__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6128__A2 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8950__A2 (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8922__A2 (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__I (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9045__A2 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9033__A3 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7974__A2 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6132__A2 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8850__B1 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7372__A2 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__I (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6130__I (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8200__B2 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7751__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__A2 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__I (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9032__A2 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7847__A2 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7843__A2 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6132__C (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8234__C (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__A2 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__C (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6134__I (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8930__A2 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7921__I (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7600__A1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__A2 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8997__A2 (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__A2 (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7866__A2 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__A2 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__B (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7658__I (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7445__I (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7025__I (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__I (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7392__B (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7337__B (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7174__B (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__B (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7949__I (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7943__I (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6360__I (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__I (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9050__B (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9047__B (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9031__B (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__A1 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8625__A1 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__I (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__A1 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6199__A1 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8922__B (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6198__A1 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9006__B (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8970__A1 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8518__A2 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__A2 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8924__A1 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8507__A1 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6996__A1 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__A1 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8850__B2 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7786__A3 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6983__I (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6152__A2 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6155__A2 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7055__I (.I(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__A1 (.I(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__A2 (.I(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7861__I (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6928__A1 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A1 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__B (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8157__C (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8106__I (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7647__I (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__C (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8513__A4 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6198__A3 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8580__A2 (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__I (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7005__A1 (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__A2 (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7769__A1 (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7063__A1 (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__B (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8779__A1 (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7076__A1 (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6191__I (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__A1 (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7182__I (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__A1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6932__A2 (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__A2 (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8520__A3 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__A2 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__A2 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__I (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__A1 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__A1 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__A1 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8932__A2 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7982__B (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7110__A2 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__I (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8006__C (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7777__I (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A2 (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__A2 (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7979__A3 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7978__A1 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__A3 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__A1 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__I (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__A1 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__A1 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7083__A2 (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__B2 (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7032__A1 (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6176__A1 (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7296__A4 (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6937__A3 (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__A3 (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6176__A2 (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7037__I (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__B (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8927__A4 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7006__A2 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6942__A2 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__A4 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8150__C (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8144__A1 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7219__A1 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__I (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7768__A1 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7733__A1 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6996__A2 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__A1 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7977__A2 (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__A2 (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9035__A3 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8507__B (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6280__A1 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__A1 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7922__A4 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__A2 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8512__A1 (.I(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__B1 (.I(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7730__B (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__A2 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__B (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6189__A2 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8963__A4 (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7879__A2 (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7035__B (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A3 (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7966__A1 (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7643__A1 (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7002__I (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6192__A1 (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7072__A1 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6940__A1 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6347__I (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6192__A2 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8929__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7721__B2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7602__I (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__A1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8990__A1 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8927__A3 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__A2 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__C (.I(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6361__A1 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__A2 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__A3 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6199__A2 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8505__A1 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7000__A2 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__I (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8925__A1 (.I(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7729__A1 (.I(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6918__A1 (.I(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6202__I (.I(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7357__I (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7237__I (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7166__I (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6203__I (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7789__A1 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7690__A1 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__B1 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6286__A1 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9028__B (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8539__A1 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__A1 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__A1 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__A2 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__A2 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__A4 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__A1 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8939__B (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__A3 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__B1 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__B2 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8938__I (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A1 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6219__B (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__B2 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__A2 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__B2 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6286__A2 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8516__A1 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7984__A1 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__A1 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6227__I (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8850__A1 (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__A1 (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__I (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__I (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8921__A1 (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7721__A1 (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7008__I (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__A1 (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8544__C (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8535__I (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6290__I (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__I (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8648__A1 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8598__B (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8562__B (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__A1 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8500__A1 (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__A2 (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8614__A1 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8595__A1 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8559__A1 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6233__A1 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8538__B (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8498__I (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__A2 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6235__I (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8997__C (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8628__A1 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8594__C (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6251__A1 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7988__A2 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__B (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__A3 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6237__I (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9015__A2 (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7884__A2 (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7878__A2 (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6243__A2 (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7985__A1 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7085__A1 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7038__A1 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6239__A1 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9006__A2 (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8996__A3 (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6243__A3 (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8257__A1 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7510__A2 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__I (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__A2 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__A1 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__A2 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__A2 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6251__A2 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8560__B (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8500__B (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6253__I (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6251__B (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__C (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9000__A2 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8887__A1 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8631__A1 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6255__A4 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__A3 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8427__A2 (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8193__A2 (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7116__I (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__I (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8292__A1 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8093__A1 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8004__A1 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__I (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8302__A1 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7324__A1 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__I (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6262__A1 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8616__A2 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8615__B (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8501__C (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6262__A2 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8630__A2 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8578__A2 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8502__A2 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__A1 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7152__A1 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7132__A1 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7121__A2 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__I (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8326__B2 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7205__A2 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6393__I (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6272__A1 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8978__A1 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7197__A1 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7190__A1 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6272__A2 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8114__A1 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8103__A1 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7254__A1 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__I (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9006__A1 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7245__A1 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__I (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6272__A3 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8155__A1 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__B2 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6307__A2 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__I (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8156__A1 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8150__A1 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7307__A1 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6271__I (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7329__B2 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7302__A1 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6959__I (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6272__A4 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7379__A1 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7355__A1 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7349__A1 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__A1 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8269__A1 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7481__B2 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7464__A1 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__I (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8630__A1 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7457__A1 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6417__I (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__A3 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__A4 (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__A1 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8935__A1 (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8531__I (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7180__A1 (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__A1 (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7808__A2 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__A2 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__A2 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__A3 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6283__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__A3 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8854__A1 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7508__A2 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7113__I (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6289__I (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7936__A1 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7789__B2 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7616__A1 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6346__A1 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8577__C (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7747__A1 (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__B1 (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__A1 (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8945__C (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8629__A1 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8598__A1 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__A1 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8921__A4 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8645__A1 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8508__A2 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__A1 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8326__C (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8062__C (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7824__I (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__A1 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8997__A1 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8944__B (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6339__A1 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6338__A3 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__C (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__A2 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8229__A1 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7405__I (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__I (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__A2 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8309__A1 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8208__A1 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8205__A1 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__A1 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9039__B (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8626__A1 (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__B2 (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8233__A1 (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7436__A1 (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6969__I (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__B1 (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8572__A1 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6307__A1 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8242__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8210__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8074__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6307__C1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__B2 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6317__A2 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8297__A1 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7672__A2 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7458__A1 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__I (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7512__A1 (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7469__A2 (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6322__B1 (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__C2 (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__A1 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7532__A1 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7514__A1 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__C2 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6330__A1 (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9005__A1 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8610__A1 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__B2 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__A1 (.I(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6322__A1 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8930__A1 (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__A1 (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__A1 (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__I (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__A1 (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__A1 (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7299__A1 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7298__B (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6954__I (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__B1 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__A2 (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8428__A1 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8092__A2 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__A1 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__A2 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8642__A1 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6338__A1 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8470__A2 (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8448__A2 (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7223__I (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6337__I (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8361__A1 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8255__A1 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A1 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6338__A2 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__A2 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8981__C (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8962__A1 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7840__A2 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__A2 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__A2 (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__C (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6358__A1 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8920__A1 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8503__C (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7899__A1 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__A1 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7896__A1 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7795__A2 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7787__A1 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__I (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7878__A1 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7850__A1 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7844__A2 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__C (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__A2 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8945__A2 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8892__A1 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8649__A1 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__A1 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8433__B2 (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7814__A2 (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7020__I (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6355__I (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8405__B2 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8386__B2 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7819__A2 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__C (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8651__A1 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__C (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7013__C (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6361__C (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6368__I (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__I (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__A2 (.I(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__A2 (.I(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__A2 (.I(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__A2 (.I(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__A2 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__A2 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__A2 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__A2 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6375__A2 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__A2 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__A2 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__A2 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7738__A1 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__A3 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8018__A2 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7862__A2 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7807__A1 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__A1 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7940__A2 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7938__A3 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6923__B (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A2 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7887__I (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6925__A2 (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__A2 (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6933__A1 (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__I (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7643__A2 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__A2 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7140__I (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6388__I (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7738__A2 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7213__A2 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6942__A1 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__A2 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__A2 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6391__I (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8991__A1 (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8989__A1 (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8502__A1 (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__A1 (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7052__A2 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7018__I (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A2 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7071__A1 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__B (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__A1 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__I (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6933__A2 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6399__I (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7283__C (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7005__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__B1 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__I (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7689__B (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7332__I (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7226__C (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6401__I (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8632__A2 (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8546__A2 (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7754__A1 (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__A2 (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8977__A1 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8545__A1 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7819__A1 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6406__A1 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8006__A1 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7957__A1 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6922__A1 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__A1 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8974__A1 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8951__A1 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8563__A1 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6411__A1 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8919__A2 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__I (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8920__A2 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8918__A2 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8917__A2 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__A2 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9033__A1 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7843__A1 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__I0 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__A1 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7975__A2 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7974__A1 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7601__A1 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6421__A1 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8392__I (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7233__I (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__A1 (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__A1 (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__A2 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__I (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__A2 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9035__A2 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9015__A1 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8784__A1 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__A1 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6591__A2 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6560__A2 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__I (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6497__A2 (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__A2 (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6443__A2 (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__A2 (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8790__B2 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__A1 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__A3 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__B1 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6876__A1 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__A1 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6443__B2 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__B2 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__A2 (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A2 (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6444__A2 (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__A2 (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__A1 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__A1 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__A1 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__A2 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6470__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6450__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__A1 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__A2 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__A2 (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__A2 (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__A1 (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__A1 (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6491__A1 (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__A2 (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6544__A1 (.I(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__B2 (.I(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__I (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__A1 (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__A1 (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__A1 (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8807__A1 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6496__A2 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6751__A2 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6750__A1 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6706__A1 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__A1 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__A2 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6509__A2 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6708__A2 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6577__B1 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__B1 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__B1 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6555__A2 (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__A2 (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__A3 (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8811__B2 (.I(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__B1 (.I(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__A1 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__A1 (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6699__A1 (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__A2 (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__I (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__A2 (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__A2 (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__A1 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6548__A1 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6747__A1 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6547__A3 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8814__B2 (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__B1 (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6749__I (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__A2 (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6696__A2 (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6573__A2 (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6812__A2 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__A1 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__A2 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__A3 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6686__A2 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6685__A2 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6588__A3 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__I (.I(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8818__B2 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__B1 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6605__I (.I(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6604__I (.I(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6595__I (.I(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6594__I (.I(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6612__A2 (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6610__A2 (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6608__A2 (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6606__A2 (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6620__I (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6615__I (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6626__A2 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6624__A2 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6622__A2 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6619__A2 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6627__A2 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6625__A2 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6623__A2 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6621__A2 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8742__A1 (.I(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8656__A1 (.I(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6888__A1 (.I(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6655__A1 (.I(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6667__I (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6666__I (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__I (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6652__I (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6663__A2 (.I(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6660__A2 (.I(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6657__A2 (.I(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6654__A2 (.I(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8744__A1 (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8658__A1 (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6890__A1 (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6658__A1 (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8746__A1 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8660__A1 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6892__A1 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6661__A1 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8748__A1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8662__A1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6894__A1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6664__A1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6677__A2 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6674__A2 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6671__A2 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6668__A2 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8754__A1 (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8668__A1 (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6900__A1 (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6672__A1 (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8756__A1 (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8670__A1 (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6902__A1 (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6675__A1 (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8758__A1 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8672__A1 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6904__A1 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6678__A1 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6678__B (.I(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6795__B1 (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6762__B1 (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6725__B1 (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6683__B1 (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6822__A1 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6793__A1 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__A1 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__A1 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6727__A1 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__A1 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8826__A1 (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__A2 (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6768__A3 (.I(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__B (.I(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6738__A1 (.I(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6833__A1 (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6812__A3 (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6811__A1 (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__A2 (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__A3 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6785__A1 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__A2 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8829__A1 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__A2 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6826__A2 (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6807__A2 (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6858__A2 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__I (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6835__A2 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6809__A2 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8835__A1 (.I(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6822__A2 (.I(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__B1 (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__A1 (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6873__A1 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6860__A3 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6858__A3 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6836__A1 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__B2 (.I(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__A2 (.I(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6878__I (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6868__A2 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__A2 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__A2 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6882__A2 (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6868__B1 (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__B1 (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__B1 (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8643__A2 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6872__A2 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6860__A2 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__A2 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6871__A2 (.I(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6865__A3 (.I(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8842__A1 (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__A2 (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8845__A1 (.I(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6876__A2 (.I(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8849__A1 (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6883__B1 (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6896__I (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6895__I (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6886__I (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6885__I (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6893__A2 (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6891__A2 (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6889__A2 (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6887__A2 (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__A2 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__A2 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__A2 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6897__A2 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8921__A2 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7814__A1 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7156__A1 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__A1 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7296__A1 (.I(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6937__A1 (.I(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__A1 (.I(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6910__A1 (.I(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7982__A2 (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7162__I (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6938__A1 (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__A1 (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7296__A3 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6937__A2 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__A2 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__A2 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7199__I (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6910__A2 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8505__A2 (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7729__A2 (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6911__A2 (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7436__B (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7149__I (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7075__A1 (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6912__I (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7669__B2 (.I(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__C (.I(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7245__B (.I(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6918__A2 (.I(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7129__I (.I(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6999__I (.I(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6915__A1 (.I(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8196__B1 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8059__A2 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6990__I (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6917__A2 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__A2 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7146__I (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6917__A3 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7795__A3 (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7081__B (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7075__A2 (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6918__A3 (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7669__A1 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7308__C (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7254__C (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__A3 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8933__A1 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7402__I (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7009__I (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6922__A2 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7909__I (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__A1 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6923__A2 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__B2 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7761__B (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__A2 (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6926__I (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8059__B (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7987__B2 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7857__I (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6932__A1 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8967__A3 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__A1 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__A2 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6928__A2 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7992__A1 (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7983__A1 (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6993__A3 (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6932__A3 (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8426__A1 (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8185__A1 (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7763__A3 (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6932__B1 (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7914__A2 (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7763__A2 (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7761__A1 (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6931__A2 (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8521__B (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7760__A2 (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__A3 (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7073__A2 (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6943__A3 (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8430__B (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8197__A1 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7743__I (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6936__A2 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6942__A3 (.I(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7642__A1 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7525__A1 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7317__B2 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6940__A2 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8851__A1 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6940__B (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6943__A4 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__S (.I(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6962__I (.I(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6948__I (.I(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6944__I (.I(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8335__A1 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7606__A1 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7539__I (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6946__I (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8000__A1 (.I(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7603__A1 (.I(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7538__A1 (.I(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6947__I (.I(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8326__A1 (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7605__A1 (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7566__B2 (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6949__A1 (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6981__A2 (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6957__A2 (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__A2 (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6949__A2 (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7605__B (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7603__A2 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7589__A1 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__A1 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7827__A1 (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7276__A1 (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7261__A2 (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6958__A1 (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8382__A1 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8379__A1 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8101__A1 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6956__I (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8398__A1 (.I(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7648__B2 (.I(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7632__A1 (.I(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6957__A1 (.I(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8917__A1 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8578__A1 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7831__A1 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6963__I0 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8401__A1 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8150__B2 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7669__C (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6961__I (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8399__A1 (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7678__B2 (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7670__A1 (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6963__I1 (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8919__A1 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8599__A1 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7835__A1 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6967__I0 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8429__A1 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7704__A1 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7702__A1 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6967__I1 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8616__A1 (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7840__A1 (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7404__A1 (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__A1 (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8453__A1 (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8232__A1 (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7798__A1 (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6971__A1 (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8472__A1 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8258__A1 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7801__A1 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__I1 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8289__A1 (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8230__A2 (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8057__A1 (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6977__I (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7598__I (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7516__A1 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7413__A2 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6978__I (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7934__A1 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7847__A1 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7689__A2 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6981__A1 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8292__B2 (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7873__B2 (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7713__B2 (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__A1 (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7907__A2 (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7906__A1 (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7868__A2 (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6989__A1 (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7983__B (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7088__A1 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7015__I (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6986__A1 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8983__A2 (.I(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8982__B (.I(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7003__A2 (.I(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6986__A2 (.I(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8971__A3 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8050__I (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7901__I (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__A2 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8934__B2 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6988__I (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8989__A2 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8977__A2 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8974__A2 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6989__A2 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__B1 (.I(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8292__B1 (.I(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8150__B1 (.I(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8101__A2 (.I(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6991__I (.I(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8925__A2 (.I(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8326__B1 (.I(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7906__A2 (.I(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__B2 (.I(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9035__A1 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7946__A1 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7014__I (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6994__A1 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7936__A3 (.I(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7876__B (.I(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6994__A2 (.I(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6997__A1 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8507__A2 (.I(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__A1 (.I(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__A1 (.I(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6996__A3 (.I(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7747__B (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6997__A2 (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__A1 (.I(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8196__A2 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7136__I (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7031__I (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7000__A1 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8934__A2 (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8486__I (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7001__I (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8623__B1 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7086__A1 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7006__A3 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7869__I (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7372__A1 (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__A1 (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7003__A1 (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8281__I (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7005__A3 (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8852__A1 (.I(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__A2 (.I(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7013__A2 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7012__C (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9011__A1 (.I(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9004__A1 (.I(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7872__A1 (.I(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7012__A1 (.I(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8430__A1 (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8054__B (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7141__A1 (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7010__I (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8402__B (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8377__A1 (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7940__A1 (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7012__A2 (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7063__A2 (.I(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7012__B (.I(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7013__B (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7929__I (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7853__A1 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7797__C (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7022__A1 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8961__B (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7939__I (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7508__A1 (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7017__I (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7897__A1 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7788__B2 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7655__B2 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7022__A2 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7073__A1 (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7056__A2 (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__A3 (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7019__I (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7871__B1 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7789__C (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7035__A2 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7022__A3 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8955__C (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7835__A2 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7831__A2 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__A2 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__A2 (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7023__A2 (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8619__B (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7855__I (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7853__A2 (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7026__I (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9040__A1 (.I(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8987__A1 (.I(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7851__A1 (.I(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7046__A1 (.I(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7062__A1 (.I(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7028__I (.I(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7797__A1 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7067__A2 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7065__A1 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__A1 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8935__A2 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8513__A3 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7924__I (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__A2 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8382__A2 (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8257__A2 (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7479__I (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7032__A2 (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__B1 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7773__A1 (.I(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7734__A1 (.I(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7044__A1 (.I(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__A2 (.I(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8584__A1 (.I(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7747__C (.I(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__A2 (.I(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7035__A1 (.I(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8342__I (.I(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8282__A1 (.I(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__A2 (.I(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8964__B (.I(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7104__I (.I(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7076__A2 (.I(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7038__A2 (.I(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8436__B2 (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8203__B2 (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8088__I (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__A3 (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7986__A1 (.I(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__A1 (.I(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8963__A2 (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__A1 (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8935__A3 (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7051__A2 (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7991__A1 (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7739__A1 (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__A2 (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7850__A2 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7805__A1 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7097__A1 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7058__A2 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7878__B (.I(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7058__A3 (.I(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8512__A2 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7805__A2 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7058__A4 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7991__A2 (.I(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7739__A2 (.I(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7059__A2 (.I(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7936__A2 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7893__A2 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7751__A2 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7072__A2 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8523__A1 (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7062__A2 (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7990__A1 (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7064__A2 (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7740__A1 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7072__B (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8924__A2 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7067__A1 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7766__I (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7069__I (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8569__I (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8494__I (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7730__A2 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7070__A2 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7087__A1 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8516__A4 (.I(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7082__A2 (.I(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8504__A1 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7994__A1 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7923__C (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7082__A3 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7760__A1 (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7736__A1 (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7178__A1 (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7081__A1 (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7882__A1 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7178__A2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7160__A2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7080__A1 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7931__A2 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7904__A2 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7882__A2 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7080__A2 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7894__B (.I(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7890__A2 (.I(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7736__A2 (.I(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7081__A2 (.I(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7994__A2 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7797__B (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7082__A4 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7989__B (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7769__A2 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7086__A3 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9015__C (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8504__B (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7850__B (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7085__B (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7741__A1 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7087__A2 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7100__A1 (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8964__A2 (.I(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7758__A1 (.I(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7737__A3 (.I(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7099__A1 (.I(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8617__A2 (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__A1 (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8011__A2 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8010__A1 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7094__A2 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8009__S (.I(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7094__B (.I(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8323__S (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8144__A2 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7859__A2 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7095__A2 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8235__A1 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8096__I (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8063__I (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7099__A2 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9034__A4 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9014__A2 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7097__A2 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7993__A2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7099__B (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7173__I (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7101__I (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7724__A2 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7692__A2 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7659__A2 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7103__I (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7447__A1 (.I(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7393__A1 (.I(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7338__A1 (.I(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7175__A1 (.I(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__B (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7286__A1 (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7170__I (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7105__I (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7801__A2 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7798__A2 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7442__A1 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7172__A1 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8009__I1 (.I(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7205__A1 (.I(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7121__A1 (.I(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7107__I (.I(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8023__A1 (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8018__A1 (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7172__B2 (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7114__A1 (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7680__I (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7109__I (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8160__B2 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8069__A1 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7144__I (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7112__A1 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8192__I (.I(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7771__I (.I(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7111__I (.I(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8403__A1 (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8359__A1 (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8327__A1 (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7112__A2 (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7715__A2 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7592__A2 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7500__A2 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7114__A2 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9010__A1 (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8946__C (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7526__A1 (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7114__B (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8380__A2 (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7727__A1 (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7520__A1 (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__I (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7496__B2 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7484__A1 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7383__A1 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7118__I (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7654__A1 (.I(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7574__A1 (.I(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7509__A1 (.I(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7126__A2 (.I(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7323__A2 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7282__A1 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__A1 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7120__I (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7874__A1 (.I(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7485__A2 (.I(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7384__A2 (.I(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__A1 (.I(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8004__A2 (.I(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__B2 (.I(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__A2 (.I(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7856__I (.I(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7781__I (.I(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7780__I (.I(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__A2 (.I(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7414__C (.I(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7125__I (.I(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7600__A2 (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7485__B (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7384__B (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7126__C (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7938__A1 (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7591__A1 (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__A1 (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7137__A1 (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8510__A1 (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8424__A2 (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7778__A1 (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7130__I (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8472__A2 (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8453__A2 (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8292__A2 (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7132__A2 (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8001__A1 (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__A2 (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7174__A1 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__A1 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7139__A1 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7138__A1 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8060__A2 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8054__A2 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7712__A2 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7135__I (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7903__I (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7875__A2 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7868__A1 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7139__A2 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8150__A2 (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8016__A1 (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7327__I (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7137__A2 (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7566__A2 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7270__I (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7212__A2 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7138__A2 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8965__A2 (.I(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7915__I (.I(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__B (.I(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7141__A2 (.I(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7566__C (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7328__B (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7142__I (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7481__C (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7376__B (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7277__B (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__C (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8387__A1 (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7788__A1 (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7655__A2 (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7145__B (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7438__A1 (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7363__A2 (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__I (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7709__A1 (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7554__A1 (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7198__B (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7167__A1 (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7629__A1 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7521__C (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7185__I (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7150__I (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7457__A2 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7308__A1 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7307__A2 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7155__A1 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7968__I (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7873__B1 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7705__A1 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7158__I (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8587__A1 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8488__A1 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7547__A1 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7159__B2 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7167__A2 (.I(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7708__A1 (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7264__I (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7161__I (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7418__A1 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7362__I (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7296__A2 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__A1 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7874__B (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7671__C (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7472__A1 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__B1 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7167__B (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8638__B (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8489__B (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7710__C (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7167__C (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7168__B (.I(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8649__A2 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8564__A2 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8525__A2 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7171__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7488__B (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7390__B (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7229__A1 (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7171__A2 (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7175__A2 (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7530__A1 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7392__A2 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7337__A2 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7174__A2 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7725__A1 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7693__A1 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7289__A1 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7235__A1 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8058__A1 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8048__A1 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7230__A1 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7226__A1 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8177__A2 (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7726__A2 (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7179__I (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7926__A2 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7527__I (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7335__I (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7180__A2 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7723__A2 (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7528__A2 (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7287__A2 (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7230__A2 (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8622__B (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7615__C (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7525__C (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7183__I (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7642__B (.I(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7565__B (.I(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7478__C (.I(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__A1 (.I(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7705__B2 (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7625__A1 (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7604__A1 (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7190__B (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7463__A1 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7437__A1 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7245__A2 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7189__A1 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7198__A1 (.I(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7516__A2 (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7455__B (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7254__A2 (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7192__I (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8621__A1 (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8604__A1 (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7355__C (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7197__C (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7198__A2 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__A2 (.I(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7634__A1 (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7614__B2 (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7439__A1 (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7207__A1 (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7232__A1 (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7224__A1 (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7212__A1 (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7201__A1 (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7211__A2 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7207__A2 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7552__I (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7524__C (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7263__A1 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7206__A1 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7207__B (.I(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__A3 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8599__C (.I(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8563__C (.I(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8545__C (.I(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7227__A2 (.I(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9016__B (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8019__A1 (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7867__A2 (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7213__A1 (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7783__A1 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7404__A2 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7377__I (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7212__B1 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7213__A3 (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8060__B1 (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7374__I (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7215__I (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8234__A1 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8151__A1 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7758__A2 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7216__A2 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7417__A2 (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7318__A2 (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7283__A2 (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7226__A2 (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8470__A3 (.I(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8056__I (.I(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__A2 (.I(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__A1 (.I(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7574__C (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7324__C (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7219__A2 (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7688__A1 (.I(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7653__B (.I(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7508__A3 (.I(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7226__B1 (.I(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8057__A2 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__A2 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8381__A1 (.I(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7572__I (.I(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7281__A2 (.I(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7224__A2 (.I(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7227__B2 (.I(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__B (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7529__A2 (.I(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7448__I (.I(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7288__A2 (.I(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7232__A2 (.I(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8484__I (.I(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8086__I (.I(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7792__I (.I(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7234__I (.I(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7756__C (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7530__C (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7289__C (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7235__C (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8649__B2 (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8630__B (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7441__A2 (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__A2 (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8587__B (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8533__B (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7440__C (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7269__A1 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8110__A1 (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7247__A1 (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7246__A1 (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7239__A1 (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__B1 (.I(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7300__A1 (.I(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7244__A1 (.I(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7243__A1 (.I(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7351__B1 (.I(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7305__A1 (.I(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7253__A1 (.I(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7252__A1 (.I(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7351__B2 (.I(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7305__A2 (.I(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7251__A1 (.I(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7254__B (.I(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7256__A2 (.I(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7269__A2 (.I(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7524__A1 (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7476__A1 (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7369__B2 (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7268__A1 (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7288__A1 (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7281__A1 (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7277__A1 (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7267__A1 (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7275__A2 (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7268__A2 (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__B (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7648__A2 (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7481__A2 (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7376__A2 (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7277__A2 (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7983__A2 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7272__I (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7987__B1 (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7496__B1 (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7326__I (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7276__A2 (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8335__A2 (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8225__A2 (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7378__I (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7274__I (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8226__A1 (.I(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7862__A3 (.I(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7714__A1 (.I(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7275__A1 (.I(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__A2 (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8093__A2 (.I(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7282__A2 (.I(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8142__A1 (.I(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7312__A1 (.I(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7311__A1 (.I(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7291__I (.I(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8146__A1 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8143__B (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7359__A1 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7336__A1 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7489__A2 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7443__A2 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7391__A2 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7336__A2 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7328__A2 (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7295__A2 (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8504__A2 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7522__I (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7438__B (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7310__A1 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__A2 (.I(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7308__A2 (.I(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7309__A3 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__B2 (.I(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8149__A2 (.I(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7324__A2 (.I(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7678__A2 (.I(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7590__A2 (.I(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7496__A2 (.I(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7329__A2 (.I(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7917__B1 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7864__B2 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7678__B1 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7329__B1 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8333__A1 (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8301__A1 (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8269__A2 (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7328__A1 (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7329__C (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8407__A1 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8094__A1 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7875__A1 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7331__B (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8580__B1 (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8564__B1 (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7441__B1 (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7333__B (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7336__B1 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7657__B2 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7617__B2 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7579__B2 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7336__B2 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8261__A2 (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7420__A1 (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7358__A1 (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7340__I (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8227__A1 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8180__A1 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7411__A1 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7341__I (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8193__A1 (.I(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8183__A1 (.I(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7391__A1 (.I(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7389__A1 (.I(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7633__A1 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7615__A1 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7478__A1 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7371__A1 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7351__A1 (.I(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7350__A1 (.I(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__A1 (.I(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7344__A1 (.I(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7434__A3 (.I(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7346__A2 (.I(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7348__A2 (.I(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7371__A2 (.I(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8606__A1 (.I(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8582__B (.I(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8551__B (.I(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7370__A1 (.I(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7466__A1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7382__A1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7364__A1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7361__A1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7466__A2 (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7364__A2 (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7361__A2 (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7965__A2 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7961__A1 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7960__A1 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7363__A1 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7392__A1 (.I(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7384__A1 (.I(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7376__A1 (.I(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7368__A1 (.I(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7398__A2 (.I(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7368__A2 (.I(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7379__B1 (.I(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7369__B1 (.I(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7370__A2 (.I(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7390__A1 (.I(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8449__B2 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8434__B2 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8201__B2 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7373__I (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8466__A3 (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8365__B2 (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7386__I (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7375__A1 (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8293__A1 (.I(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7681__A2 (.I(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7649__A2 (.I(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7375__A2 (.I(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7577__A2 (.I(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7487__A2 (.I(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7389__A2 (.I(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7648__B1 (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7566__B1 (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7481__B1 (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7379__A2 (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8302__A2 (.I(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7679__A1 (.I(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7499__A1 (.I(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7379__B2 (.I(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7568__A2 (.I(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7482__A2 (.I(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7410__A2 (.I(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7382__A2 (.I(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8194__A2 (.I(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7383__A2 (.I(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8305__B2 (.I(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7575__B (.I(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7487__B2 (.I(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7389__B2 (.I(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9002__B (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8177__A1 (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7796__A1 (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7388__I (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8942__A1 (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7898__C (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7487__C (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7389__C (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7391__B (.I(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8286__A2 (.I(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7468__A1 (.I(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7408__A1 (.I(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7395__I (.I(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8230__A1 (.I(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8228__A1 (.I(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7443__A1 (.I(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7441__A1 (.I(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8157__A1 (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8115__A1 (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8055__A1 (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7400__A1 (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7494__A3 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7474__A2 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7399__A2 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7439__A2 (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7400__A2 (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7474__A1 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7446__A1 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7413__A1 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__A1 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8922__A1 (.I(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8383__B (.I(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8259__B (.I(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__C (.I(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7415__A1 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8400__S (.I(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8290__A2 (.I(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8058__A2 (.I(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7406__I (.I(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8325__A2 (.I(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8324__A1 (.I(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7507__A2 (.I(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7414__A1 (.I(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8266__A1 (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8265__A1 (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7423__A1 (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7408__A2 (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8229__A2 (.I(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7414__A2 (.I(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8329__A1 (.I(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8095__A1 (.I(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7745__A2 (.I(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7417__B2 (.I(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7710__A1 (.I(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7676__A1 (.I(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7440__A1 (.I(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7568__A3 (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7482__A3 (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7422__A1 (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7433__A1 (.I(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7432__A1 (.I(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7426__A1 (.I(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7425__A1 (.I(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7794__I (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7607__A1 (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7450__I (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7431__C (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7438__A2 (.I(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7437__A2 (.I(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7438__A3 (.I(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7439__B (.I(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7441__C (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7443__B (.I(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7660__A1 (.I(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7619__A1 (.I(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7581__A1 (.I(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7491__A1 (.I(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8262__A1 (.I(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7510__A1 (.I(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7489__A1 (.I(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7487__A1 (.I(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8605__A1 (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8581__A1 (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8550__A1 (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7465__A1 (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8298__A1 (.I(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7673__A2 (.I(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7637__B (.I(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7452__A1 (.I(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7463__A2 (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7478__A2 (.I(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7558__A1 (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7482__B (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7471__A3 (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7470__A2 (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7490__A1 (.I(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7485__A1 (.I(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7481__A1 (.I(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7475__A1 (.I(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7480__A2 (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7476__A2 (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7488__A1 (.I(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8326__A2 (.I(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8270__A1 (.I(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7646__A1 (.I(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7480__A1 (.I(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7504__A2 (.I(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7483__A2 (.I(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8255__A2 (.I(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7484__A2 (.I(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7489__B (.I(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8321__A1 (.I(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8295__A1 (.I(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7528__A1 (.I(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7500__A1 (.I(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7529__A1 (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7507__A1 (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7496__A1 (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7495__A1 (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7524__A2 (.I(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7499__A2 (.I(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8967__A4 (.I(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7498__I (.I(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7714__C (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7679__C (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7591__C (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7499__C (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7556__A2 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7511__A1 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7506__A1 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7558__C (.I(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7505__A1 (.I(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7526__B (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7519__A3 (.I(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7738__B2 (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7670__C (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7523__B (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7524__B (.I(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7526__C (.I(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7790__A1 (.I(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7723__B2 (.I(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7691__B2 (.I(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7528__B2 (.I(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7691__A2 (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7657__A2 (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7617__A2 (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7579__A2 (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8334__A1 (.I(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7609__A1 (.I(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__A1 (.I(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7554__A2 (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7580__A1 (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7573__A1 (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7566__A1 (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7551__A1 (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7567__A2 (.I(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7553__A2 (.I(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7969__A3 (.I(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7934__A3 (.I(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7883__A1 (.I(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7553__B (.I(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7578__A1 (.I(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7570__A1 (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7569__B (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7563__A1 (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7561__A1 (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7568__A4 (.I(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7559__A2 (.I(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7558__A2 (.I(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7558__B (.I(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7560__A2 (.I(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7709__C (.I(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7634__C (.I(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7614__A1 (.I(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7564__A1 (.I(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7567__B (.I(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7575__A1 (.I(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7570__A3 (.I(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7569__A2 (.I(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7716__A1 (.I(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7651__A1 (.I(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7596__A2 (.I(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7571__A1 (.I(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8324__A2 (.I(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7574__A2 (.I(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8466__A2 (.I(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7687__A1 (.I(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7653__A2 (.I(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7573__A2 (.I(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8617__C (.I(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7683__B (.I(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7655__C (.I(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7577__B (.I(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7578__B2 (.I(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7579__B1 (.I(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7581__B (.I(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8370__A1 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7637__A1 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7617__A1 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7592__A1 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8401__A2 (.I(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8103__A2 (.I(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7589__A2 (.I(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7584__I (.I(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8607__A1 (.I(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8588__A1 (.I(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8485__I (.I(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7588__A1 (.I(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7618__A1 (.I(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7599__A1 (.I(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7590__A1 (.I(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7587__A1 (.I(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7614__B1 (.I(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7588__A2 (.I(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7592__B1 (.I(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8362__A1 (.I(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7591__A2 (.I(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8361__A2 (.I(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7601__A2 (.I(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7785__A1 (.I(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7720__A2 (.I(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7719__A1 (.I(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7599__A2 (.I(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7720__B (.I(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7601__C (.I(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8650__A2 (.I(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8589__A2 (.I(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7942__A1 (.I(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7616__B2 (.I(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8378__A1 (.I(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8353__A1 (.I(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8059__A1 (.I(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7609__B (.I(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7615__A2 (.I(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7614__A2 (.I(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7615__B (.I(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7616__C (.I(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7617__B1 (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8422__A2 (.I(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8380__A1 (.I(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7673__A1 (.I(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7621__I (.I(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8410__A1 (.I(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8375__A1 (.I(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7657__A1 (.I(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7655__A1 (.I(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7665__A2 (.I(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7624__A2 (.I(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7632__A2 (.I(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8424__A3 (.I(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7701__A4 (.I(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7627__I (.I(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7670__A2 (.I(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7632__B (.I(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7634__B (.I(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7656__A1 (.I(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8434__C (.I(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8201__C (.I(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7644__I (.I(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8449__C (.I(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8365__C (.I(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7682__B2 (.I(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7645__I (.I(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8406__A1 (.I(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8305__C (.I(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7870__A1 (.I(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7650__A1 (.I(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7649__B1 (.I(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8475__A1 (.I(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8447__A1 (.I(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8158__A1 (.I(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7648__C (.I(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7649__B2 (.I(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8381__A2 (.I(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7654__A2 (.I(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7947__B (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7724__B (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7692__B (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7659__B (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8417__A1 (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8411__A1 (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7691__A1 (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7681__A1 (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7692__A1 (.I(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7689__A1 (.I(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7678__A1 (.I(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7666__A1 (.I(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7679__A2 (.I(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7671__A2 (.I(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7671__B (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7677__A1 (.I(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7683__A1 (.I(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8272__B2 (.I(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8238__B2 (.I(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8023__B1 (.I(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7682__A2 (.I(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7690__B (.I(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8400__I1 (.I(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7687__A2 (.I(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8443__A1 (.I(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8427__A1 (.I(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7723__A1 (.I(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7715__A1 (.I(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7710__A2 (.I(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7709__A2 (.I(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7714__A2 (.I(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7708__A2 (.I(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7722__A1 (.I(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8446__A1 (.I(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8425__A1 (.I(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7712__A1 (.I(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7713__B1 (.I(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7715__B (.I(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8428__A2 (.I(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7719__A2 (.I(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7720__C (.I(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7723__B1 (.I(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7954__I (.I(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7941__C (.I(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7738__B1 (.I(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7729__B1 (.I(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7957__B (.I(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7728__I (.I(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8852__A2 (.I(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7734__A2 (.I(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8928__A3 (.I(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7986__A3 (.I(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7734__A3 (.I(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7957__C (.I(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7933__A3 (.I(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7732__A2 (.I(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8851__A2 (.I(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8505__B (.I(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7733__B (.I(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7740__A2 (.I(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7738__C (.I(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7742__A2 (.I(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7756__A1 (.I(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7755__A2 (.I(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8377__A2 (.I(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8236__B2 (.I(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8152__A1 (.I(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7744__I (.I(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8404__B2 (.I(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8271__C (.I(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7911__A2 (.I(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7746__A1 (.I(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7747__A2 (.I(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7746__A2 (.I(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8481__A1 (.I(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8344__A1 (.I(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8131__C (.I(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7753__A1 (.I(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7934__A2 (.I(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7933__A2 (.I(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7874__A2 (.I(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__A2 (.I(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7883__C (.I(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__C (.I(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8972__A1 (.I(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7765__A2 (.I(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7992__A2 (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7762__A2 (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7894__A2 (.I(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7762__A3 (.I(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7994__B (.I(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7765__B (.I(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7774__A3 (.I(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8626__A2 (.I(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8590__A2 (.I(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8572__A2 (.I(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7768__A2 (.I(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8476__C (.I(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8473__C (.I(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8453__C (.I(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7772__A1 (.I(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8384__B2 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8260__A1 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8103__B1 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7772__A2 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7774__A4 (.I(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7776__A2 (.I(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7905__A1 (.I(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7786__A2 (.I(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7784__A2 (.I(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7779__A2 (.I(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7982__C (.I(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7940__A3 (.I(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7782__A2 (.I(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7779__A3 (.I(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8435__A1 (.I(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8202__A1 (.I(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8020__A1 (.I(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7785__A2 (.I(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8159__A1 (.I(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8067__B (.I(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7894__A1 (.I(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7784__A3 (.I(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7992__A3 (.I(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7783__A2 (.I(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8047__C (.I(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7803__C (.I(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7800__C (.I(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7793__C (.I(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8586__A1 (.I(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8549__I (.I(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8532__A1 (.I(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7795__A1 (.I(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7803__A1 (.I(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7802__A2 (.I(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7800__A1 (.I(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7799__A2 (.I(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8921__A3 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8339__A1 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7881__I (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7809__A1 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9016__A1 (.I(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7880__A1 (.I(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7871__A1 (.I(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7808__B2 (.I(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7821__I (.I(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7811__I (.I(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7810__I (.I(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8959__A1 (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8950__A1 (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7839__A2 (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7813__A2 (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8943__A2 (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7815__A2 (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8548__A1 (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7820__A1 (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7979__A2 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7969__A1 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7832__A2 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7820__A2 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9030__A1 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7822__I0 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9034__A1 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8992__A2 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7836__A2 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7827__A2 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8944__A2 (.I(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8363__B (.I(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8263__A1 (.I(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7826__A2 (.I(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9010__A2 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7828__I0 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8585__A1 (.I(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7832__A1 (.I(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9048__A1 (.I(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9024__A1 (.I(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7832__B (.I(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9049__A1 (.I(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9025__A1 (.I(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7833__A2 (.I(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9042__A1 (.I(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9019__A1 (.I(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7836__B (.I(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9046__A1 (.I(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9021__A1 (.I(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7837__A2 (.I(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8997__B (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7841__I0 (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9039__A1 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7846__A2 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7846__A3 (.I(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7848__I0 (.I(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7981__A2 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7972__A2 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7900__A2 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7880__A2 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8417__B (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8346__B (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8137__B (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7879__A1 (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8477__A1 (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8376__B (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8117__A1 (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7871__A2 (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8065__A1 (.I(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7912__I (.I(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7891__I (.I(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7858__I (.I(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8062__A1 (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8019__C (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7864__A1 (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7863__B (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8364__A1 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8264__A1 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7895__A2 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7864__A2 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7930__A4 (.I(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7865__I (.I(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7863__A1 (.I(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7862__A1 (.I(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9018__A1 (.I(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7914__A1 (.I(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7876__A1 (.I(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7867__A1 (.I(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7896__A2 (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7867__B (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7870__B1 (.I(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8957__B2 (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8918__A1 (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7917__C (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7870__B2 (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7882__A3 (.I(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7877__A1 (.I(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7883__B (.I(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7877__A2 (.I(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7878__C (.I(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7879__A4 (.I(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9045__A1 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9033__A2 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9020__A1 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7884__A1 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7884__B (.I(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8983__C (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8616__C (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8502__C (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7886__I (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8503__A1 (.I(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8341__A1 (.I(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8119__A1 (.I(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7898__A1 (.I(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8412__A1 (.I(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8358__B (.I(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8329__C (.I(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7895__A1 (.I(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8220__A1 (.I(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8065__B (.I(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8001__B (.I(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7889__I (.I(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8355__A1 (.I(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8354__A1 (.I(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8271__A1 (.I(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7890__A1 (.I(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8968__A1 (.I(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8104__C (.I(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8066__A1 (.I(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7892__I (.I(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8456__A1 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8303__B2 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8116__C (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7893__A1 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7900__B1 (.I(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8366__B1 (.I(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8120__I (.I(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8042__A2 (.I(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7902__I (.I(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8958__A1 (.I(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8440__A1 (.I(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8215__A1 (.I(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7908__A1 (.I(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8636__A1 (.I(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8623__A1 (.I(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7911__A1 (.I(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7907__A1 (.I(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8328__A1 (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8151__B2 (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7940__B (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7911__A3 (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7927__A1 (.I(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7923__A2 (.I(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7914__C (.I(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7911__A4 (.I(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8433__A1 (.I(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8200__A1 (.I(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8158__C (.I(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7913__I (.I(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8376__A1 (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8338__C (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7917__B2 (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7914__B (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8409__A1 (.I(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8236__C (.I(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8095__C (.I(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7916__I (.I(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8340__C (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8304__A1 (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8273__A1 (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7917__A2 (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8459__A1 (.I(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8391__A1 (.I(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8284__A1 (.I(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7920__B (.I(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9044__A1 (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8340__A1 (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7977__B (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7922__A2 (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7923__B (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8366__A2 (.I(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8204__I (.I(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8041__I (.I(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7925__I (.I(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8457__A2 (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8415__A2 (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8131__B2 (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7926__A1 (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7941__B (.I(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7935__A1 (.I(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7937__A1 (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7937__A2 (.I(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8984__A1 (.I(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8617__A1 (.I(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8415__B2 (.I(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7941__A1 (.I(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9027__C (.I(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9023__C (.I(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7965__B (.I(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7944__C (.I(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8441__C (.I(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8317__C (.I(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8216__C (.I(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7950__I (.I(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8483__A1 (.I(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8461__A1 (.I(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8371__A1 (.I(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7953__A1 (.I(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7971__A2 (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7969__B (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7964__A1 (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7963__A2 (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8238__A1 (.I(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8160__A1 (.I(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8023__A2 (.I(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7956__I (.I(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8467__A1 (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8387__B2 (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8272__A1 (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7957__A2 (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7964__A2 (.I(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7961__A2 (.I(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7960__A2 (.I(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7963__B (.I(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8434__A1 (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8201__A1 (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8068__A1 (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7967__I (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8449__A1 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8365__A1 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8305__A1 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7971__A1 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8638__A1 (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8533__A1 (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8489__A1 (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7969__A2 (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7971__B1 (.I(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7978__B2 (.I(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7985__A2 (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8972__A2 (.I(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7984__A2 (.I(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7990__A4 (.I(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8135__A1 (.I(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7996__A1 (.I(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7995__A1 (.I(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7994__C (.I(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8135__A2 (.I(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7996__A2 (.I(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8440__B (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8316__B (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8215__B (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7998__I (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8250__A2 (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8175__A2 (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8087__A2 (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8047__A2 (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8249__A1 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8174__A1 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8085__A1 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8046__A2 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8015__A1 (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8360__A2 (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8254__A2 (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8149__A1 (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8003__A2 (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8023__B2 (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8006__A2 (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8097__A2 (.I(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8064__A2 (.I(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8008__A2 (.I(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8969__A2 (.I(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8967__A2 (.I(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8220__A2 (.I(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8014__I (.I(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8385__B2 (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8355__C (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8263__C (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8015__B (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8020__A2 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8019__A2 (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8238__C (.I(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8160__C (.I(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8069__C (.I(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8022__I (.I(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8467__C (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8387__C (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8272__C (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8023__C (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8044__A1 (.I(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8244__A1 (.I(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8161__I (.I(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8079__B1 (.I(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8027__I (.I(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8310__A1 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8209__A1 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8206__A1 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8029__A1 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8311__B2 (.I(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8308__A2 (.I(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8207__A2 (.I(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8032__B2 (.I(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8308__B1 (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8274__B1 (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8170__A2 (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8039__A2 (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8240__A1 (.I(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8126__B2 (.I(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8122__B2 (.I(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8037__B2 (.I(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8491__A2 (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8042__B1 (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8247__B2 (.I(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8172__B2 (.I(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8082__B2 (.I(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8042__B2 (.I(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8480__A1 (.I(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8458__A1 (.I(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8283__A1 (.I(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8044__B (.I(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8176__I (.I(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8174__C (.I(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8085__C (.I(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8046__C (.I(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8085__A2 (.I(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8068__A2 (.I(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8066__B2 (.I(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8051__A2 (.I(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8313__A1 (.I(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8247__A1 (.I(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8141__A1 (.I(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8051__A1 (.I(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8055__A2 (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8362__A2 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8055__B (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8062__A2 (.I(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8431__B2 (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8291__A1 (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8100__A1 (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8061__A1 (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8069__A2 (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8061__A2 (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8067__A1 (.I(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8433__A2 (.I(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8263__B2 (.I(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8200__A2 (.I(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8066__A2 (.I(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8066__A3 (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8303__A1 (.I(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8237__A1 (.I(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8182__I (.I(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8066__B1 (.I(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8082__A2 (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8309__B2 (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8208__B2 (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8205__B2 (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8071__B2 (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8311__C (.I(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8210__C (.I(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8128__B (.I(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8074__C (.I(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8207__B1 (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8128__A2 (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8124__A2 (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8080__A2 (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8079__A1 (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8243__A1 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8240__B2 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8126__A1 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8078__A1 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8541__A2 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8082__B1 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8390__C (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8248__B (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8173__B (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8084__B (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8285__C (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8250__C (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8175__C (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8087__C (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8416__A1 (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8345__A1 (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8316__A1 (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8134__A1 (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8134__A2 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8116__A2 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8103__B2 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8131__A2 (.I(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8104__A2 (.I(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8095__A2 (.I(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8100__A2 (.I(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8094__A2 (.I(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8474__A1 (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8376__A2 (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8358__A1 (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8105__A1 (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8143__A2 (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8142__A3 (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8098__A2 (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8105__A2 (.I(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8473__A1 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8455__A1 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8147__A1 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8104__A1 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8104__B2 (.I(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8446__C (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8269__B (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8115__C (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8107__I (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8476__A1 (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8338__A1 (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8337__A1 (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8116__A1 (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8115__A2 (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8258__A2 (.I(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8233__A2 (.I(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8156__A2 (.I(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8114__A2 (.I(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8116__B (.I(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8479__A1 (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8457__B1 (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8390__B1 (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8131__A1 (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8557__A2 (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8131__B1 (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8134__B2 (.I(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8391__C (.I(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8284__C (.I(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8249__C (.I(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8133__I (.I(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8441__A2 (.I(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8416__C (.I(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8345__C (.I(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8134__C (.I(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8481__C (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8368__I (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8136__I (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8417__A2 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8370__A2 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8346__A2 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8137__A2 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8217__A3 (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8179__A2 (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8146__A2 (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8140__A2 (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8174__A2 (.I(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8158__A2 (.I(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8141__A2 (.I(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8261__A3 (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8227__A2 (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8183__A2 (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8145__A1 (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8455__B2 (.I(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8412__A2 (.I(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8296__B2 (.I(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8145__B (.I(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8151__C (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8157__A2 (.I(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8158__B (.I(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8172__A2 (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8307__A1 (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8278__A1 (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8169__B1 (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8164__A1 (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8540__A1 (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8277__B2 (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8168__B2 (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8163__B2 (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8952__A2 (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8279__B2 (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8274__A2 (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8166__B2 (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8574__A2 (.I(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8172__B1 (.I(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8394__A2 (.I(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8317__A2 (.I(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8285__A2 (.I(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8216__A2 (.I(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8414__B (.I(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8178__I (.I(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8439__A1 (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8369__A1 (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8315__A1 (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8214__A1 (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8180__A2 (.I(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8198__A2 (.I(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8181__I (.I(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8215__A2 (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8214__A2 (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8203__A2 (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8201__A2 (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8436__A1 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8405__A1 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8386__A1 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8203__A1 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8200__A3 (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8223__A2 (.I(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8191__A2 (.I(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8190__A2 (.I(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8199__A2 (.I(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8472__B1 (.I(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8452__A1 (.I(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8431__A1 (.I(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8198__A1 (.I(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8201__B1 (.I(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8198__B1 (.I(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8453__B1 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8256__I (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8231__A1 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8198__B2 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8197__A2 (.I(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8198__C (.I(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8199__B (.I(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8200__B1 (.I(_3364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8437__A2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8390__A2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8313__B2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8212__A1 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8592__A2 (.I(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8212__A2 (.I(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8213__A2 (.I(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8249__A2 (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8247__A2 (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8234__A2 (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8238__A2 (.I(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8237__A2 (.I(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8302__B (.I(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8236__A1 (.I(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8226__A2 (.I(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8236__A2 (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8238__B1 (.I(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8231__A2 (.I(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8446__B (.I(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8233__B (.I(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8234__B (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8237__B (.I(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8611__A2 (.I(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8247__B1 (.I(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8284__A2 (.I(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8282__A2 (.I(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8272__A2 (.I(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8264__A2 (.I(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8272__B1 (.I(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8260__B1 (.I(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8403__B2 (.I(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8384__A1 (.I(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8362__B2 (.I(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8260__B2 (.I(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8259__A1 (.I(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8475__A2 (.I(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8259__A2 (.I(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8260__C (.I(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8263__B1 (.I(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8270__A2 (.I(_3431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8271__B (.I(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8276__A2 (.I(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8627__A2 (.I(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8282__B1 (.I(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8957__A2 (.I(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8478__A2 (.I(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8343__A2 (.I(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8282__B2 (.I(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8318__A2 (.I(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8287__A2 (.I(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8316__A2 (.I(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8313__A2 (.I(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8305__A2 (.I(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8288__I (.I(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8290__B (.I(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8293__C (.I(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8356__A3 (.I(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8321__A2 (.I(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8295__A2 (.I(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8296__B1 (.I(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8302__C (.I(_3463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8303__C (.I(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8640__A2 (.I(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8313__B1 (.I(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8349__A2 (.I(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8348__A3 (.I(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8319__A2 (.I(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8345__A2 (.I(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8343__B2 (.I(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8340__A2 (.I(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8338__A2 (.I(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8322__A2 (.I(_3482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8339__A2 (.I(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8328__A2 (.I(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8328__B (.I(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8341__A2 (.I(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8378__A2 (.I(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8353__A2 (.I(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8336__A2 (.I(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8337__A2 (.I(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8338__B (.I(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8993__B (.I(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8990__A2 (.I(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8414__A1 (.I(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8343__B1 (.I(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8366__B2 (.I(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8359__A2 (.I(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8352__I (.I(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8369__A2 (.I(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8365__A2 (.I(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8364__A2 (.I(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8355__A2 (.I(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8354__A2 (.I(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8365__B1 (.I(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8362__B1 (.I(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8367__B (.I(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8482__A2 (.I(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8460__A2 (.I(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8459__C (.I(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8369__C (.I(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8384__B1 (.I(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8373__I (.I(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8376__A3 (.I(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8404__A1 (.I(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8385__A1 (.I(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8385__A2 (.I(_3538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8387__A2 (.I(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8384__A2 (.I(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8384__C (.I(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8386__B1 (.I(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8890__I (.I(_3551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8869__I (.I(_3551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8602__I (.I(_3551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8393__I (.I(_3551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8585__C (.I(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8566__C (.I(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8548__C (.I(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8394__C (.I(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8416__A2 (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8414__A2 (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8408__A2 (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8405__A2 (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8404__A2 (.I(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8403__C (.I(_3560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8405__B1 (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8415__B1 (.I(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8420__A2 (.I(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8440__A2 (.I(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8439__A2 (.I(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8436__A2 (.I(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8434__A2 (.I(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8450__A2 (.I(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8423__A2 (.I(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8446__A2 (.I(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8425__A2 (.I(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8432__A1 (.I(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8434__B1 (.I(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8431__B1 (.I(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8430__A2 (.I(_3586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8431__C (.I(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8438__A2 (.I(_3594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8457__A1 (.I(_3598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8458__A2 (.I(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8457__B2 (.I(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8455__A2 (.I(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8447__A2 (.I(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8447__B (.I(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8473__A2 (.I(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8467__A2 (.I(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8479__C (.I(_3633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9013__A1 (.I(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8976__A1 (.I(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8949__A1 (.I(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8528__A1 (.I(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8527__A1 (.I(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8499__A1 (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8553__I (.I(_3646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8538__A1 (.I(_3646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8508__A1 (.I(_3646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8493__I (.I(_3646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8926__A2 (.I(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8593__B (.I(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8557__C (.I(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8497__A1 (.I(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8641__A2 (.I(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8609__A2 (.I(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8554__A2 (.I(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8496__A2 (.I(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8496__B (.I(_3649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8499__A2 (.I(_3651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8500__A2 (.I(_3653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8527__A2 (.I(_3657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8515__A3 (.I(_3659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8508__A4 (.I(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8514__A2 (.I(_3662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8510__B2 (.I(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8511__A2 (.I(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8514__A3 (.I(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8523__A3 (.I(_3669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8580__C (.I(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8529__I (.I(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8526__I (.I(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8524__I (.I(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8649__C (.I(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8600__A1 (.I(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8546__B (.I(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8525__B (.I(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8528__A2 (.I(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8619__A1 (.I(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8603__A2 (.I(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8565__A1 (.I(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8530__I (.I(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8631__A2 (.I(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8618__A2 (.I(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8601__A2 (.I(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8547__A2 (.I(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8547__B (.I(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8615__A1 (.I(_3689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8567__I (.I(_3689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8544__A1 (.I(_3689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8543__A1 (.I(_3689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8866__A1 (.I(_3690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8576__A2 (.I(_3690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8564__A1 (.I(_3690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8544__A2 (.I(_3690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8542__B2 (.I(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8543__A2 (.I(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8546__C (.I(_3698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8548__B (.I(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8565__A2 (.I(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8591__A2 (.I(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8556__A2 (.I(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8558__B (.I(_3709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8560__A1 (.I(_3710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8646__A1 (.I(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8628__C (.I(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8576__C (.I(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8562__A1 (.I(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8564__C (.I(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8566__B (.I(_3717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9000__A1 (.I(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8999__A1 (.I(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8946__A1 (.I(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8577__A1 (.I(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8965__A1 (.I(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8627__C (.I(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8612__A1 (.I(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8574__C (.I(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8576__B1 (.I(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8577__B (.I(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8584__C (.I(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8585__B (.I(_3735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8601__B (.I(_3738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8594__B (.I(_3743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8596__A1 (.I(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8883__A1 (.I(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8628__A2 (.I(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8618__A1 (.I(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8598__A2 (.I(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8600__A3 (.I(_3749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8865__C (.I(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8861__C (.I(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8634__C (.I(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8603__C (.I(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8618__B (.I(_3756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8614__A2 (.I(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8998__A1 (.I(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8614__B (.I(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8618__C (.I(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8620__B (.I(_3768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8628__B2 (.I(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8629__B (.I(_3776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8632__C (.I(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8645__A2 (.I(_3791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8646__C (.I(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8650__C (.I(_3796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8664__I (.I(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8663__I (.I(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8654__I (.I(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8653__I (.I(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8661__A2 (.I(_3800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8659__A2 (.I(_3800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8657__A2 (.I(_3800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8655__A2 (.I(_3800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8671__A2 (.I(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8669__A2 (.I(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8667__A2 (.I(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8665__A2 (.I(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8764__A1 (.I(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8724__A1 (.I(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8705__A1 (.I(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8680__A1 (.I(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8682__I (.I(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8676__I (.I(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8698__A2 (.I(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8695__A2 (.I(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8678__I (.I(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8677__I (.I(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8690__A2 (.I(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8687__A2 (.I(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8684__A2 (.I(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8680__A2 (.I(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8699__A2 (.I(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8696__A2 (.I(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8693__A2 (.I(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8679__A2 (.I(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8767__A1 (.I(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8727__A1 (.I(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8708__A1 (.I(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8684__A1 (.I(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8692__A2 (.I(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8689__A2 (.I(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8686__A2 (.I(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8683__A2 (.I(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8769__A1 (.I(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8729__A1 (.I(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8710__A1 (.I(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8687__A1 (.I(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8771__A1 (.I(_3823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8731__A1 (.I(_3823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8712__A1 (.I(_3823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8690__A1 (.I(_3823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8773__A1 (.I(_3825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8733__A1 (.I(_3825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8714__A1 (.I(_3825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8693__A1 (.I(_3825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8775__A1 (.I(_3827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8735__A1 (.I(_3827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8716__A1 (.I(_3827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8696__A1 (.I(_3827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8777__A1 (.I(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8737__A1 (.I(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8718__A1 (.I(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8699__A1 (.I(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8706__I (.I(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8701__I (.I(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8712__A2 (.I(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8710__A2 (.I(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8708__A2 (.I(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8705__A2 (.I(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8718__A2 (.I(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8716__A2 (.I(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8714__A2 (.I(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8704__A2 (.I(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8713__A2 (.I(_3836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8711__A2 (.I(_3836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8709__A2 (.I(_3836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8707__A2 (.I(_3836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8725__I (.I(_3843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8720__I (.I(_3843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8731__A2 (.I(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8729__A2 (.I(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8727__A2 (.I(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8724__A2 (.I(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8732__A2 (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8730__A2 (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8728__A2 (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8726__A2 (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8750__I (.I(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8749__I (.I(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8740__I (.I(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8739__I (.I(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8765__I (.I(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8760__I (.I(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8771__A2 (.I(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8769__A2 (.I(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8767__A2 (.I(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8764__A2 (.I(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8777__A2 (.I(_3871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8775__A2 (.I(_3871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8773__A2 (.I(_3871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8763__A2 (.I(_3871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8772__A2 (.I(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8770__A2 (.I(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8768__A2 (.I(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8766__A2 (.I(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8822__A1 (.I(_3880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8806__A1 (.I(_3880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8786__A1 (.I(_3880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8820__A1 (.I(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8784__A2 (.I(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8808__A2 (.I(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8799__A2 (.I(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8795__A2 (.I(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8790__A2 (.I(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8825__I (.I(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8818__B1 (.I(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8798__I (.I(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8789__I (.I(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8845__A2 (.I(_3891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8842__A2 (.I(_3891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8795__B1 (.I(_3891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8790__B1 (.I(_3891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8815__A2 (.I(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8812__A2 (.I(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8809__A2 (.I(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8792__I (.I(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8804__A2 (.I(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8800__A2 (.I(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8796__A2 (.I(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8793__A2 (.I(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8849__A2 (.I(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8840__A2 (.I(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8807__A2 (.I(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8849__B2 (.I(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8819__A1 (.I(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8835__A2 (.I(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8832__A2 (.I(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8829__A2 (.I(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8826__A2 (.I(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8847__I (.I(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8844__A2 (.I(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8841__A2 (.I(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8839__A2 (.I(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8848__A2 (.I(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8844__B1 (.I(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8841__B1 (.I(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8839__B1 (.I(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8880__I (.I(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8875__I (.I(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8859__I (.I(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8853__I (.I(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8877__I (.I(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8876__I (.I(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8856__I (.I(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8855__I (.I(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8861__A2 (.I(_3944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8865__A2 (.I(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8870__A2 (.I(_3951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8874__A2 (.I(_3955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8895__A1 (.I(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8891__A1 (.I(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8886__A1 (.I(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8882__A1 (.I(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8882__A2 (.I(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8886__A2 (.I(_3965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8891__A2 (.I(_3968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9005__C (.I(_3970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8995__C (.I(_3970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8895__C (.I(_3970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8891__C (.I(_3970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8895__A2 (.I(_3972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8908__I (.I(_3974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8907__I (.I(_3974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8898__I (.I(_3974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8897__I (.I(_3974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8906__A1 (.I(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8904__A1 (.I(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8902__A1 (.I(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8900__A1 (.I(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8905__A2 (.I(_3976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8903__A2 (.I(_3976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8901__A2 (.I(_3976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8899__A2 (.I(_3976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9007__A1 (.I(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8936__A1 (.I(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8928__A2 (.I(_3993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9007__A2 (.I(_3996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8936__A2 (.I(_3996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9006__C (.I(_3997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8931__A1 (.I(_3997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9007__A3 (.I(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8936__A4 (.I(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8996__B (.I(_4004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8937__A2 (.I(_4004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8948__A2 (.I(_4005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8947__A3 (.I(_4005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8942__A3 (.I(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8973__A1 (.I(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8966__A3 (.I(_4030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8970__A2 (.I(_4034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8973__A3 (.I(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8989__B (.I(_4040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8977__B (.I(_4040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8974__B (.I(_4040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8981__B (.I(_4046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8987__A2 (.I(_4052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8993__A2 (.I(_4057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9005__A2 (.I(_4060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9004__B (.I(_4060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8998__A2 (.I(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9003__A2 (.I(_4065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9002__A2 (.I(_4065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9004__C (.I(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9012__A2 (.I(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9011__C (.I(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9011__A2 (.I(_4071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9017__A1 (.I(_4077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9036__A1 (.I(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9017__A2 (.I(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9029__I (.I(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9028__A2 (.I(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9024__A2 (.I(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9019__A2 (.I(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9030__A3 (.I(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9025__A2 (.I(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9021__A2 (.I(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9048__A2 (.I(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9042__A2 (.I(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9039__A2 (.I(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9038__B (.I(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9040__A2 (.I(_4098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9049__A2 (.I(_4103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9046__A2 (.I(_4103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__S (.I(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__S (.I(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5649__S (.I(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__I (.I(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__S (.I(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__S1 (.I(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__I (.I(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__I (.I(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__S1 (.I(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__S1 (.I(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__S (.I(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__I (.I(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A1 (.I(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__I (.I(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__A1 (.I(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__A1 (.I(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8778__B (.I(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6138__I (.I(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__A2 (.I(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__A2 (.I(_4117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__I (.I(_4117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__A2 (.I(_4117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__A2 (.I(_4117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8780__A1 (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__A1 (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__A1 (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A1 (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__I (.I(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__A2 (.I(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A2 (.I(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4544__A1 (.I(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__A2 (.I(_4123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__I (.I(_4123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__A3 (.I(_4123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A2 (.I(_4123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__A1 (.I(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6158__I (.I(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4544__A2 (.I(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__A2 (.I(_4125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__I (.I(_4125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__I (.I(_4125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7061__A1 (.I(_4126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__A2 (.I(_4126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__I (.I(_4126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A2 (.I(_4126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__A1 (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__A3 (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__A1 (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__I (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__I (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__I (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__A2 (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__S (.I(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A2 (.I(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__I (.I(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__I (.I(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__A2 (.I(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__A2 (.I(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__A1 (.I(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__I (.I(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__I (.I(_4132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__A1 (.I(_4132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__A1 (.I(_4132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__I (.I(_4132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7096__A1 (.I(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__A1 (.I(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__A1 (.I(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__A1 (.I(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__A1 (.I(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__A2 (.I(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__I (.I(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__A1 (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__I (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A2 (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__A1 (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__A1 (.I(_4136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__A1 (.I(_4136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__I (.I(_4136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__I (.I(_4136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__I (.I(_4137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__I (.I(_4137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__A1 (.I(_4137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__A2 (.I(_4137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8521__A1 (.I(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__A1 (.I(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__A1 (.I(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__A1 (.I(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6150__I (.I(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__A1 (.I(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__A3 (.I(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__A2 (.I(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4712__I (.I(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A2 (.I(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7096__A2 (.I(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__A2 (.I(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__A1 (.I(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__A2 (.I(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__S0 (.I(_4146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__S0 (.I(_4146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A1 (.I(_4146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__I (.I(_4146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__A1 (.I(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6243__A1 (.I(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A1 (.I(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__A1 (.I(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6294__A1 (.I(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__A2 (.I(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__A1 (.I(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__A3 (.I(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__A2 (.I(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4759__A1 (.I(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__A1 (.I(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__I (.I(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__A1 (.I(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__I (.I(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__A1 (.I(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__A1 (.I(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4710__A1 (.I(_4155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__A1 (.I(_4155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A1 (.I(_4155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__A1 (.I(_4155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__A2 (.I(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__A1 (.I(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__A2 (.I(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7049__A2 (.I(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6062__I (.I(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__A3 (.I(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__A1 (.I(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__I (.I(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__I (.I(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__C (.I(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__A2 (.I(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__I (.I(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__A1 (.I(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__A2 (.I(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__I (.I(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__I (.I(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__A1 (.I(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__I (.I(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__A2 (.I(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9035__A4 (.I(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6156__A2 (.I(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__A2 (.I(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__A2 (.I(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8497__B2 (.I(_4169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7047__A2 (.I(_4169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__A1 (.I(_4169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__I (.I(_4169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7733__A2 (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5888__A1 (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__A1 (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__A2 (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__A1 (.I(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6060__A1 (.I(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__A1 (.I(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__A1 (.I(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A2 (.I(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__I (.I(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__A2 (.I(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__A1 (.I(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__S0 (.I(_4173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__I (.I(_4173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__A1 (.I(_4173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__A1 (.I(_4173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A2 (.I(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__I (.I(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__A2 (.I(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__A2 (.I(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__A2 (.I(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__I (.I(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__A2 (.I(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__A2 (.I(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__A2 (.I(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__I (.I(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__A1 (.I(_4177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__A2 (.I(_4177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__I (.I(_4177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__A2 (.I(_4177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8779__A2 (.I(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__A1 (.I(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__I (.I(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__A2 (.I(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__A2 (.I(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__I (.I(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__I (.I(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__A2 (.I(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__A2 (.I(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__I (.I(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A2 (.I(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8012__A1 (.I(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8011__C (.I(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7094__A1 (.I(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__A1 (.I(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__A1 (.I(_4184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__A1 (.I(_4184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4621__A1 (.I(_4184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__I (.I(_4184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__A1 (.I(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6152__A1 (.I(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__A1 (.I(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__A1 (.I(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__A1 (.I(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__A1 (.I(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__I (.I(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__A2 (.I(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7955__I (.I(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__A2 (.I(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7944__A2 (.I(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7931__B (.I(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__A1 (.I(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A1 (.I(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6913__A1 (.I(_4190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__A4 (.I(_4190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A1 (.I(_4190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A3 (.I(_4190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__I (.I(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__A2 (.I(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A1 (.I(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7011__A1 (.I(_4193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6157__I (.I(_4193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__A1 (.I(_4193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__A2 (.I(_4193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7214__A2 (.I(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6921__I (.I(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6915__A2 (.I(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A1 (.I(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6422__A1 (.I(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__A2 (.I(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4710__A2 (.I(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__A1 (.I(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8007__A2 (.I(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__I (.I(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__I (.I(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__A1 (.I(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__A1 (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__A3 (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__I (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__A2 (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7066__A2 (.I(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__A2 (.I(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__A2 (.I(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6995__I (.I(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__A2 (.I(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__A1 (.I(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__A2 (.I(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__I (.I(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__A3 (.I(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4621__A2 (.I(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8927__A1 (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7006__A1 (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__A2 (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A2 (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8518__C (.I(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__A2 (.I(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__B (.I(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__A1 (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__A2 (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7095__A1 (.I(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__I (.I(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__A1 (.I(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__A1 (.I(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__A1 (.I(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__I (.I(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A1 (.I(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__I (.I(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6925__A1 (.I(_4210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__A1 (.I(_4210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__A1 (.I(_4210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__A1 (.I(_4210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5563__A1 (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__B2 (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__A1 (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__A2 (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__A1 (.I(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__A1 (.I(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__A1 (.I(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__A2 (.I(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A1 (.I(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__I (.I(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__A1 (.I(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A1 (.I(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A3 (.I(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__A2 (.I(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__I (.I(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A4 (.I(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6110__I (.I(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A2 (.I(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A1 (.I(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__A3 (.I(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__I (.I(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__I (.I(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7058__A1 (.I(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__I (.I(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A1 (.I(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__A2 (.I(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__B2 (.I(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5570__B (.I(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A1 (.I(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7098__A1 (.I(_4224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7047__A1 (.I(_4224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__A2 (.I(_4224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__A1 (.I(_4224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__A2 (.I(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__A2 (.I(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6173__I (.I(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A1 (.I(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7068__A1 (.I(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__I (.I(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__A1 (.I(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__I (.I(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7066__A1 (.I(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__A2 (.I(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__A1 (.I(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A2 (.I(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7809__A2 (.I(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__A2 (.I(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A3 (.I(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__A2 (.I(_4229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__A3 (.I(_4229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__I (.I(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__I (.I(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A2 (.I(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6156__A1 (.I(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__A2 (.I(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__I (.I(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__I (.I(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__A1 (.I(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__A1 (.I(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__I (.I(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8932__A1 (.I(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8517__B (.I(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7083__A1 (.I(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__A1 (.I(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6906__I (.I(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__I (.I(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__A1 (.I(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A1 (.I(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7763__A1 (.I(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__A2 (.I(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__A1 (.I(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A1 (.I(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7930__A1 (.I(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5617__A1 (.I(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__A1 (.I(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__A3 (.I(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6908__I (.I(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__A2 (.I(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__I (.I(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A2 (.I(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7430__I (.I(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A1 (.I(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8854__A2 (.I(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__A2 (.I(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__A2 (.I(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7153__I (.I(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A2 (.I(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5880__A1 (.I(_4247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__I (.I(_4247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8517__A2 (.I(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7628__A1 (.I(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5950__A1 (.I(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__A3 (.I(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7011__A2 (.I(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__A1 (.I(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__A1 (.I(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__I (.I(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8511__A1 (.I(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7056__A1 (.I(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6238__I (.I(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__A1 (.I(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__A3 (.I(_4252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__I (.I(_4252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__A1 (.I(_4252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__A1 (.I(_4252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5603__I (.I(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__I (.I(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8190__B (.I(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7397__I (.I(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7134__I (.I(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__A2 (.I(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8782__A1 (.I(_4257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7057__A1 (.I(_4257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__A2 (.I(_4257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__A2 (.I(_4257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__A2 (.I(_4258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__I (.I(_4258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__A1 (.I(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5460__A2 (.I(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__I (.I(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__A3 (.I(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__A2 (.I(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__A2 (.I(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__I (.I(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8510__A2 (.I(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__I (.I(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__A2 (.I(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__A4 (.I(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__A3 (.I(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__A3 (.I(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8505__C (.I(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5970__A1 (.I(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5934__A1 (.I(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__A2 (.I(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7876__A2 (.I(_4267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__A2 (.I(_4267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__A2 (.I(_4267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__I (.I(_4268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__A1 (.I(_4268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__I (.I(_4268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8779__A3 (.I(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8517__A1 (.I(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8516__A3 (.I(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__A2 (.I(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__A1 (.I(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5705__I (.I(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A1 (.I(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__A2 (.I(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7807__A2 (.I(_4271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__A1 (.I(_4271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__I (.I(_4271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__A2 (.I(_4273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__A1 (.I(_4273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__I (.I(_4273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5534__A1 (.I(_4276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__A2 (.I(_4276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__A1 (.I(_4276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__I (.I(_4276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7543__A1 (.I(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__A4 (.I(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A2 (.I(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__I (.I(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8520__A2 (.I(_4278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7297__I (.I(_4278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7243__B (.I(_4278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A2 (.I(_4278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__I (.I(_4280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__A3 (.I(_4280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__A2 (.I(_4282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__I (.I(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6142__I (.I(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__C (.I(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__C (.I(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__C (.I(_4288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A1 (.I(_4288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__A1 (.I(_4288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__A1 (.I(_4288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__B (.I(_4289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__I (.I(_4289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__I (.I(_4289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4709__I (.I(_4289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__A2 (.I(_4291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4759__A2 (.I(_4291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__I (.I(_4291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__A1 (.I(_4292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__A1 (.I(_4292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__A2 (.I(_4292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A1 (.I(_4292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__A2 (.I(_4293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A2 (.I(_4293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__A2 (.I(_4293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A2 (.I(_4293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6183__I (.I(_4294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__A3 (.I(_4294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__A3 (.I(_4294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__A2 (.I(_4294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__A1 (.I(_4295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__A3 (.I(_4295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__I (.I(_4295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A3 (.I(_4295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__C (.I(_4297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5098__I (.I(_4297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__C (.I(_4297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__I (.I(_4297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8942__A2 (.I(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5480__B2 (.I(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__B2 (.I(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__A1 (.I(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__A1 (.I(_4299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6450__A1 (.I(_4299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__I (.I(_4299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__A1 (.I(_4299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__A1 (.I(_4300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__B1 (.I(_4300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__I (.I(_4300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__B1 (.I(_4300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__A1 (.I(_4301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__S (.I(_4301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__S1 (.I(_4301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__S (.I(_4301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8052__A2 (.I(_4302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8016__A2 (.I(_4302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__B2 (.I(_4302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__A1 (.I(_4303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__A1 (.I(_4303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__I (.I(_4303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__C1 (.I(_4303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__C2 (.I(_4304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__C (.I(_4305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__I (.I(_4305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__I (.I(_4305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__I (.I(_4305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__I (.I(_4306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__A2 (.I(_4306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__A2 (.I(_4306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__A2 (.I(_4306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__A1 (.I(_4309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__A1 (.I(_4309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__A1 (.I(_4309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__I (.I(_4309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__A1 (.I(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__A1 (.I(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A1 (.I(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__I (.I(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__A1 (.I(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6154__A1 (.I(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__A1 (.I(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__A1 (.I(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8934__A1 (.I(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__A2 (.I(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__A2 (.I(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__A2 (.I(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__A1 (.I(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__A1 (.I(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__A1 (.I(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__A1 (.I(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__A1 (.I(_4315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4750__A1 (.I(_4315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__B2 (.I(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__A2 (.I(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__A2 (.I(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__I (.I(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__A1 (.I(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__I (.I(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__A1 (.I(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__A1 (.I(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__B (.I(_4319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__A1 (.I(_4319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__A2 (.I(_4319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__I (.I(_4319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7816__A1 (.I(_4322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__I0 (.I(_4322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__A1 (.I(_4322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__A1 (.I(_4322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__A3 (.I(_4324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A3 (.I(_4324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__A3 (.I(_4324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6223__A1 (.I(_4330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A2 (.I(_4330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__A2 (.I(_4330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4750__A2 (.I(_4330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__A2 (.I(_4333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__B (.I(_4333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__B (.I(_4333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__I (.I(_4333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9001__A1 (.I(_4334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__A1 (.I(_4334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__A1 (.I(_4334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__A1 (.I(_4334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8496__A1 (.I(_4335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__A1 (.I(_4335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__A2 (.I(_4335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__B (.I(_4336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__A1 (.I(_4336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__B (.I(_4336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__A1 (.I(_4336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__B2 (.I(_4338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__B2 (.I(_4338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__I (.I(_4338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A1 (.I(_4338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6156__A3 (.I(_4340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__I (.I(_4340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__A1 (.I(_4341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__A1 (.I(_4341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__A1 (.I(_4341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A2 (.I(_4341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8490__A2 (.I(_4347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6204__A1 (.I(_4347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__A1 (.I(_4347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A2 (.I(_4347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__C (.I(_4349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__I (.I(_4349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__I (.I(_4349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__I (.I(_4349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__C (.I(_4351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5432__C (.I(_4351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__C (.I(_4351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4771__I (.I(_4351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7813__A1 (.I(_4353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__B2 (.I(_4353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6244__A3 (.I(_4353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4773__I (.I(_4353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8944__A1 (.I(_4354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5920__A1 (.I(_4354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__I (.I(_4354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__A1 (.I(_4354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__A1 (.I(_4356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__I (.I(_4356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__A1 (.I(_4356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9026__A1 (.I(_4357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8570__A1 (.I(_4357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__A1 (.I(_4357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A1 (.I(_4357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6830__A1 (.I(_4358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6742__A1 (.I(_4358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6696__A1 (.I(_4358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__I (.I(_4358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6786__A1 (.I(_4359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A1 (.I(_4359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__I (.I(_4359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__A1 (.I(_4359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__A1 (.I(_4361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__A1 (.I(_4361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__A1 (.I(_4361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4781__I (.I(_4361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__I (.I(_4362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A2 (.I(_4362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5413__A1 (.I(_4362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__A1 (.I(_4362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8331__A2 (.I(_4363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8330__A2 (.I(_4363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8300__A2 (.I(_4363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__A2 (.I(_4363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__A2 (.I(_4364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4789__A2 (.I(_4364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__S0 (.I(_4366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__S0 (.I(_4366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__S0 (.I(_4366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__I (.I(_4366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__A1 (.I(_4367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__A2 (.I(_4367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__I (.I(_4367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__S0 (.I(_4367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__A2 (.I(_4368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8629__A2 (.I(_4370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__A1 (.I(_4370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__A1 (.I(_4370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A2 (.I(_4370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6231__A2 (.I(_4371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5919__A1 (.I(_4371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__A2 (.I(_4371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__A1 (.I(_4372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__A3 (.I(_4372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__A1 (.I(_4372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__A2 (.I(_4372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__I (.I(_4373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__I (.I(_4373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__I (.I(_4373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__A1 (.I(_4375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__I (.I(_4375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__S (.I(_4375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__S1 (.I(_4375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__A2 (.I(_4376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__A2 (.I(_4377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__A1 (.I(_4377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__I (.I(_4377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__A1 (.I(_4378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__A2 (.I(_4378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__A1 (.I(_4378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__A1 (.I(_4378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__A1 (.I(_4379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__I (.I(_4379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4947__I (.I(_4379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A1 (.I(_4379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8110__A2 (.I(_4380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8109__A2 (.I(_4380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8053__A2 (.I(_4380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__B2 (.I(_4380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__A3 (.I(_4381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__A2 (.I(_4381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__I (.I(_4381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__A2 (.I(_4382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__A3 (.I(_4382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__A2 (.I(_4382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__A2 (.I(_4382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__A1 (.I(_4383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__I (.I(_4383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__I (.I(_4384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__A1 (.I(_4384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A1 (.I(_4384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__A2 (.I(_4384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8781__A1 (.I(_4385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__C (.I(_4385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__I (.I(_4385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__A1 (.I(_4385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7204__A2 (.I(_4386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7187__A1 (.I(_4386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__A2 (.I(_4386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__I (.I(_4386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__A1 (.I(_4387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__A2 (.I(_4387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__I (.I(_4387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__A1 (.I(_4387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__I (.I(_4388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__A2 (.I(_4388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5599__I (.I(_4389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__A1 (.I(_4389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6122__A1 (.I(_4391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__A2 (.I(_4391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8506__A2 (.I(_4392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__I (.I(_4392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6261__I (.I(_4392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__A2 (.I(_4392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8963__A1 (.I(_4393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__A1 (.I(_4393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__A2 (.I(_4393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5910__A1 (.I(_4394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__A2 (.I(_4394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__I (.I(_4395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__I (.I(_4395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__A2 (.I(_4395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__I (.I(_4395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__B (.I(_4397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__I1 (.I(_4397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__I (.I(_4397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4817__I (.I(_4397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8946__A2 (.I(_4398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__A2 (.I(_4398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__A1 (.I(_4398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__A2 (.I(_4398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8503__A2 (.I(_4399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7090__A1 (.I(_4399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5916__B2 (.I(_4399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__A1 (.I(_4399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__B2 (.I(_4403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__A1 (.I(_4403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__A1 (.I(_4403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__A1 (.I(_4403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__A2 (.I(_4404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__I (.I(_4404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__A2 (.I(_4404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__A1 (.I(_4404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8516__A2 (.I(_4405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__I (.I(_4405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__A1 (.I(_4405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__A2 (.I(_4405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__A2 (.I(_4406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__I (.I(_4406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__A1 (.I(_4406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8850__A2 (.I(_4408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7873__A2 (.I(_4408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7750__I (.I(_4408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__A2 (.I(_4408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8568__I (.I(_4409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__A2 (.I(_4409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7208__I (.I(_4410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7034__I (.I(_4410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6154__A2 (.I(_4410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__A3 (.I(_4410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8781__A3 (.I(_4413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__I (.I(_4413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7732__A1 (.I(_4420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A2 (.I(_4420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6036__I (.I(_4420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__A1 (.I(_4420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6936__C (.I(_4421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5631__I (.I(_4421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__B (.I(_4421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__A1 (.I(_4421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__A1 (.I(_4422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__A2 (.I(_4422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__A2 (.I(_4422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7731__A2 (.I(_4425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6919__I (.I(_4425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6911__A1 (.I(_4425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__A1 (.I(_4425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7731__A1 (.I(_4427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7210__A1 (.I(_4427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6979__I (.I(_4427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__A1 (.I(_4427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__A2 (.I(_4429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__A3 (.I(_4429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8783__A3 (.I(_4430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__A1 (.I(_4430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__I (.I(_4430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4850__I (.I(_4430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__A1 (.I(_4436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__I (.I(_4436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__A1 (.I(_4436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__A2 (.I(_4436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8488__A2 (.I(_4438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7155__A2 (.I(_4438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5921__A1 (.I(_4438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__A2 (.I(_4438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9022__A1 (.I(_4442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__A1 (.I(_4442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__A1 (.I(_4442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__A1 (.I(_4442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7982__A1 (.I(_4443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7972__A1 (.I(_4443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7970__A1 (.I(_4443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__A1 (.I(_4443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7963__A1 (.I(_4444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7933__A1 (.I(_4444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7873__A1 (.I(_4444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__A2 (.I(_4444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__A1 (.I(_4445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5939__A1 (.I(_4445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__A3 (.I(_4445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8779__A4 (.I(_4446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7186__I (.I(_4446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__A2 (.I(_4446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__I (.I(_4446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7436__A2 (.I(_4447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7184__I (.I(_4447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7151__A1 (.I(_4447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__A2 (.I(_4447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__A1 (.I(_4449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__C (.I(_4449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__A1 (.I(_4449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__A1 (.I(_4450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__I (.I(_4450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__A1 (.I(_4450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__A1 (.I(_4450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7802__A1 (.I(_4451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__A1 (.I(_4451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__I (.I(_4451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__A1 (.I(_4451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7799__A1 (.I(_4452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__A2 (.I(_4452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__A2 (.I(_4452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__I (.I(_4452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__A2 (.I(_4453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__A2 (.I(_4453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__A1 (.I(_4455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__A1 (.I(_4455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7187__A2 (.I(_4458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__I (.I(_4458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8489__A2 (.I(_4459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7151__A2 (.I(_4459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__A1 (.I(_4459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__A2 (.I(_4459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8824__A1 (.I(_4463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8793__A1 (.I(_4463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__A2 (.I(_4463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8782__A2 (.I(_4464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__A1 (.I(_4464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__A1 (.I(_4464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8591__B (.I(_4465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8556__B (.I(_4465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6193__A1 (.I(_4465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__I (.I(_4465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8981__A1 (.I(_4466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8955__A1 (.I(_4466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8954__C (.I(_4466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__I (.I(_4466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8992__A3 (.I(_4467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5530__A2 (.I(_4467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__A1 (.I(_4467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__A2 (.I(_4467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8275__S (.I(_4468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__A1 (.I(_4468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__I (.I(_4468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__I (.I(_4468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8079__A2 (.I(_4471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8025__A1 (.I(_4471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__I (.I(_4471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__I (.I(_4471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5518__B2 (.I(_4473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__A2 (.I(_4473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__A2 (.I(_4473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__I (.I(_4473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__B2 (.I(_4474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__B2 (.I(_4474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__A1 (.I(_4474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__A2 (.I(_4474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8169__A2 (.I(_4475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__I (.I(_4475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__A2 (.I(_4475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__I (.I(_4475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__A2 (.I(_4476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__B2 (.I(_4476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__A2 (.I(_4476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__A1 (.I(_4476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__A1 (.I(_4477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__I (.I(_4477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__A1 (.I(_4477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__A1 (.I(_4477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8495__A1 (.I(_4478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__A1 (.I(_4478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__B2 (.I(_4478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__B2 (.I(_4478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8025__A2 (.I(_4483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__I (.I(_4483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__A2 (.I(_4483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__I (.I(_4483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__B1 (.I(_4484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__B1 (.I(_4484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__A2 (.I(_4484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__I (.I(_4484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__A2 (.I(_4485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__A2 (.I(_4485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__A2 (.I(_4485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__A2 (.I(_4485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8279__C (.I(_4488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8166__C (.I(_4488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8032__C (.I(_4488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__I (.I(_4488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__C (.I(_4489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__C (.I(_4489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__B (.I(_4489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__I (.I(_4489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8957__A1 (.I(_4490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__B (.I(_4490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__B (.I(_4490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__B (.I(_4490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8952__A1 (.I(_4494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5518__A1 (.I(_4494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__A1 (.I(_4494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__I (.I(_4494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8674__A1 (.I(_4495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6592__I (.I(_4495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__A1 (.I(_4495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__A1 (.I(_4495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8245__C (.I(_4497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8207__C (.I(_4497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8080__B (.I(_4497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__I (.I(_4497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8276__B (.I(_4498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8170__B (.I(_4498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5518__C (.I(_4498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__I (.I(_4498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8955__A2 (.I(_4499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__A1 (.I(_4499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__A1 (.I(_4499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__C (.I(_4499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8343__A1 (.I(_4501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__I1 (.I(_4501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__A3 (.I(_4501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8992__A1 (.I(_4503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__A1 (.I(_4503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__I (.I(_4503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__A1 (.I(_4503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7068__A2 (.I(_4504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__A1 (.I(_4504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8571__I (.I(_4506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__A2 (.I(_4506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__I (.I(_4506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8627__A1 (.I(_4508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8574__A1 (.I(_4508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5169__I (.I(_4508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__I (.I(_4508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__A2 (.I(_4510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__A1 (.I(_4510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__A2 (.I(_4510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__A2 (.I(_4510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7093__A1 (.I(_4512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A1 (.I(_4512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__A2 (.I(_4512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8506__A3 (.I(_4514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7070__A1 (.I(_4514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A2 (.I(_4514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__A2 (.I(_4514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9043__A1 (.I(_4515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9034__A2 (.I(_4515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__A2 (.I(_4515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8806__B (.I(_4517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__A1 (.I(_4517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__B (.I(_4517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__B (.I(_4517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__B (.I(_4519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__A2 (.I(_4522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__I (.I(_4522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__A2 (.I(_4522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7626__A2 (.I(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7608__I (.I(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7606__A2 (.I(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__I (.I(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8424__A1 (.I(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7703__A1 (.I(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7701__A1 (.I(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6960__I (.I(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8196__B2 (.I(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7711__I (.I(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__I (.I(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4854__A2 (.I(\as2650.addr_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__I (.I(\as2650.addr_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__I (.I(\as2650.addr_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__I (.I(\as2650.addr_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__A1 (.I(\as2650.addr_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__I (.I(\as2650.addr_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__I (.I(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__A1 (.I(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__A1 (.I(\as2650.alu_op[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__A1 (.I(\as2650.alu_op[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__I (.I(\as2650.alu_op[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__I (.I(\as2650.alu_op[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__A1 (.I(\as2650.alu_op[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__I (.I(\as2650.alu_op[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__A2 (.I(\as2650.alu_op[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A2 (.I(\as2650.alu_op[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__I (.I(\as2650.alu_op[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7945__I (.I(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__A2 (.I(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__A4 (.I(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__A4 (.I(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6907__I (.I(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__A1 (.I(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__A2 (.I(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__A2 (.I(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__I (.I(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__A1 (.I(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__A1 (.I(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7822__I1 (.I(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A1 (.I(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__A1 (.I(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7828__I1 (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__A1 (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__A1 (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__I (.I(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__A1 (.I(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7841__I1 (.I(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__A1 (.I(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__A1 (.I(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7845__A1 (.I(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__A1 (.I(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__A1 (.I(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7848__I1 (.I(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__A1 (.I(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__A1 (.I(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__I (.I(\as2650.idx_ctrl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__A2 (.I(\as2650.idx_ctrl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__A2 (.I(\as2650.idx_ctrl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__I (.I(\as2650.idx_ctrl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__A1 (.I(\as2650.idx_ctrl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__A1 (.I(\as2650.idx_ctrl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4578__A2 (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__I (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__A1 (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__A1 (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A3 (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__I (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9012__A1 (.I(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8554__A1 (.I(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__B2 (.I(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8139__A3 (.I(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__I (.I(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7620__I (.I(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5667__I (.I(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7696__A1 (.I(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7661__I (.I(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5679__I (.I(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8462__A2 (.I(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7699__A1 (.I(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7694__I (.I(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__I (.I(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8462__A1 (.I(\as2650.pc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8448__A1 (.I(\as2650.pc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8444__A1 (.I(\as2650.pc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__I (.I(\as2650.pc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8139__A2 (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7258__A1 (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7203__A1 (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5742__I (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8139__A1 (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__A1 (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__I (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7290__I (.I(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5760__I (.I(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7339__I (.I(\as2650.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__I (.I(\as2650.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8286__A1 (.I(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7503__A1 (.I(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__I (.I(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7501__A1 (.I(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5792__I (.I(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8348__A2 (.I(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7637__A2 (.I(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7555__A1 (.I(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__I (.I(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6323__I (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__I (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__A1 (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__A1 (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__A2 (.I(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__A2 (.I(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__I (.I(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__I (.I(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8556__A1 (.I(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A1 (.I(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__I (.I(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__I (.I(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9042__B (.I(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8591__A1 (.I(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__I (.I(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8609__A1 (.I(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__B2 (.I(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__A1 (.I(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6128__A1 (.I(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8641__A1 (.I(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7975__A1 (.I(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7973__I (.I(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__A1 (.I(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6573__A1 (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__B2 (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__A1 (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__I (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__B2 (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6519__A1 (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6467__I (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__I (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6577__B2 (.I(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6514__A1 (.I(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__A1 (.I(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__I (.I(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6542__A1 (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__I (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6576__A1 (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__I (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__A1 (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__I (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6579__A1 (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5408__I (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__A1 (.I(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__A1 (.I(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__A1 (.I(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__I (.I(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__I0 (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__I (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__I1 (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__I (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__I1 (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__I0 (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__I (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__I1 (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__I0 (.I(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__I (.I(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__I1 (.I(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__I (.I(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__I1 (.I(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__I3 (.I(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__I (.I(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5649__I1 (.I(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__I3 (.I(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__I (.I(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__I1 (.I(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__I3 (.I(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5976__I (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5674__A2 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__I3 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__I (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__I1 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__I3 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__I (.I(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__A2 (.I(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__I (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__A2 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__I3 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__I1 (.I(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__I (.I(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__I3 (.I(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__A1 (.I(\as2650.r123_2[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__I2 (.I(\as2650.r123_2[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__A1 (.I(\as2650.r123_2[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__I2 (.I(\as2650.r123_2[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6497__A1 (.I(\as2650.r123_2[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__I2 (.I(\as2650.r123_2[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__A1 (.I(\as2650.r123_2[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__A2 (.I(\as2650.r123_2[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__A1 (.I(\as2650.r123_2[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__I2 (.I(\as2650.r123_2[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__A1 (.I(\as2650.r123_2[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__I2 (.I(\as2650.r123_2[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6683__B2 (.I(\as2650.r123_2[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__I1 (.I(\as2650.r123_2[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8028__A2 (.I(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__A1 (.I(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A1 (.I(\as2650.stack[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__A2 (.I(\as2650.stack[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__A1 (.I(\as2650.stack[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__A1 (.I(\as2650.stack[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8909__A1 (.I(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8210__B1 (.I(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8911__A1 (.I(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8242__B1 (.I(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8913__A1 (.I(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8279__B1 (.I(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8915__A1 (.I(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8311__B1 (.I(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5661__A1 (.I(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__A1 (.I(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8242__A2 (.I(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6671__A1 (.I(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8279__A2 (.I(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6674__A1 (.I(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8726__A1 (.I(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__A1 (.I(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8078__B1 (.I(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6889__A1 (.I(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8243__B1 (.I(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__A1 (.I(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8306__B1 (.I(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__A1 (.I(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8243__A2 (.I(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6608__A1 (.I(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8306__A2 (.I(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6612__A1 (.I(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__A1 (.I(\as2650.stack[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__A1 (.I(\as2650.stack[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6377__A1 (.I(\as2650.stack[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__A1 (.I(\as2650.stack[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8661__A1 (.I(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8167__I (.I(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8741__A1 (.I(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8039__A1 (.I(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8772__A1 (.I(\as2650.stack[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__A1 (.I(\as2650.stack[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8776__A1 (.I(\as2650.stack[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5512__A1 (.I(\as2650.stack[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8743__A1 (.I(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8080__A1 (.I(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8745__A1 (.I(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8124__A1 (.I(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8747__A1 (.I(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8170__A1 (.I(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8751__A1 (.I(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8207__B2 (.I(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8753__A1 (.I(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8245__B2 (.I(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8757__A1 (.I(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8308__B2 (.I(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8766__A1 (.I(\as2650.stack[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__A1 (.I(\as2650.stack[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[33]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7407__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7503__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7501__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6311__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6315__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7979__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7976__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8052__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7221__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7238__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7203__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7312__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7311__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7424__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7420__A2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7409__A2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output14_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output15_I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output16_I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output18_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output19_I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8885__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output20_I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8889__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output21_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8894__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7023__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output23_I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7045__A1 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output24_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6982__I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout49_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout50_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout54_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output28_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output29_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7293__A2 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7266__A1 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7200__I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output30_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7293__A1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7265__I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout53_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output31_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output32_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7398__A1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7366__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output33_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7494__A2 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7401__I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7399__A1 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output34_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7494__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7473__I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output35_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7549__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7493__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output36_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7623__A2 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7586__A1 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7548__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7623__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7585__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout52_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output38_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output39_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7706__A1 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7664__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout51_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output40_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout46_I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout47_I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9382__I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9379__I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7791__A1 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7786__A1 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7784__A1 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7779__A1 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7755__A1 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__A1 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7745__A1 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7724__A1 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7720__A1 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7713__A1 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7707__A1 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7659__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7653__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7648__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7622__I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7337__A1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7329__A1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7322__I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7294__A1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7293__A3 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7266__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7133__I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7115__I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9164__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9299__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9301__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9297__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9300__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9161__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9298__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9160__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9163__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9162__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9165__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9296__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9128__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9166__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9303__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9304__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9208__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9242__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9302__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9210__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9206__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9204__CLK (.I(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9207__CLK (.I(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9167__CLK (.I(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9119__CLK (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9323__CLK (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9118__CLK (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9237__CLK (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9205__CLK (.I(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9328__CLK (.I(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9209__CLK (.I(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9211__CLK (.I(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9055__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9054__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9051__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9052__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9329__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9053__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9289__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9290__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9117__CLK (.I(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9106__CLK (.I(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9322__CLK (.I(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9327__CLK (.I(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9203__CLK (.I(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9182__CLK (.I(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9202__CLK (.I(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9244__CLK (.I(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9177__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9179__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9180__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9183__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9178__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9176__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9181__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9185__CLK (.I(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9311__CLK (.I(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9309__CLK (.I(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9312__CLK (.I(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9310__CLK (.I(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9223__CLK (.I(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9222__CLK (.I(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9220__CLK (.I(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9224__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9234__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9226__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9235__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9236__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9233__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9261__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9285__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9263__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9283__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9268__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9256__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9254__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9257__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9266__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9260__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9259__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9253__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9255__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9262__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9267__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9265__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9258__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9264__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9287__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9282__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9288__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9215__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9214__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9105__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9212__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9325__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9251__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9324__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9326__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9064__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9221__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9279__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9278__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9280__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9281__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9249__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9250__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9252__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9070__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9078__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9073__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9081__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9071__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9159__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9156__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9158__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9175__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9157__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9172__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9074__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9077__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9069__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9080__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9072__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9079__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9152__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9155__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9315__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9314__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9316__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9313__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9271__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9273__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9272__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9065__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9059__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9063__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9269__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9284__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9108__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9113__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9061__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9137__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9090__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9142__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9111__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9270__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9139__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9112__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9092__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9062__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9060__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9138__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9109__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9110__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9277__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9248__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9247__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9246__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9168__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9245__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9154__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9275__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9153__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9276__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9096__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9143__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9141__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9274__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9129__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9171__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9169__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9170__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9132__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9131__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9088__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9085__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9150__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9145__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9144__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9320__CLK (.I(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9136__CLK (.I(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9134__CLK (.I(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9133__CLK (.I(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9135__CLK (.I(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9334__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9332__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9330__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9333__CLK (.I(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9321__CLK (.I(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9099__CLK (.I(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9098__CLK (.I(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9097__CLK (.I(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9100__CLK (.I(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9123__CLK (.I(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9291__CLK (.I(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9122__CLK (.I(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9121__CLK (.I(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9124__CLK (.I(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9125__CLK (.I(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9294__CLK (.I(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9295__CLK (.I(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9292__CLK (.I(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_1_0_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_65_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9331__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_wb_clk_i_I (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_wb_clk_i_I (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_wb_clk_i_I (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_wb_clk_i_I (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9120__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_wb_clk_i_I (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_wb_clk_i_I (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_3_0_wb_clk_i_I (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_2_0_wb_clk_i_I (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9184__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_wb_clk_i_I (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_wb_clk_i_I (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_4_0_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_5_0_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9227__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9225__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9200__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9213__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9218__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9230__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_wb_clk_i_I (.I(clknet_opt_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_wb_clk_i_I (.I(clknet_opt_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9194__CLK (.I(clknet_opt_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_wb_clk_i_I (.I(clknet_opt_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_wb_clk_i_I (.I(clknet_opt_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1577 ();
 assign io_oeb[0] = net85;
 assign io_oeb[13] = net90;
 assign io_oeb[14] = net55;
 assign io_oeb[15] = net56;
 assign io_oeb[16] = net57;
 assign io_oeb[17] = net58;
 assign io_oeb[18] = net59;
 assign io_oeb[19] = net60;
 assign io_oeb[1] = net86;
 assign io_oeb[20] = net61;
 assign io_oeb[21] = net62;
 assign io_oeb[22] = net63;
 assign io_oeb[23] = net64;
 assign io_oeb[24] = net65;
 assign io_oeb[25] = net66;
 assign io_oeb[26] = net67;
 assign io_oeb[27] = net68;
 assign io_oeb[28] = net69;
 assign io_oeb[29] = net70;
 assign io_oeb[2] = net87;
 assign io_oeb[30] = net71;
 assign io_oeb[31] = net72;
 assign io_oeb[32] = net73;
 assign io_oeb[33] = net91;
 assign io_oeb[34] = net92;
 assign io_oeb[35] = net93;
 assign io_oeb[36] = net94;
 assign io_oeb[37] = net95;
 assign io_oeb[3] = net88;
 assign io_oeb[4] = net89;
 assign io_out[0] = net74;
 assign io_out[13] = net79;
 assign io_out[1] = net75;
 assign io_out[2] = net76;
 assign io_out[33] = net80;
 assign io_out[34] = net81;
 assign io_out[35] = net82;
 assign io_out[36] = net83;
 assign io_out[37] = net84;
 assign io_out[3] = net77;
 assign io_out[4] = net78;
endmodule

