VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO avali_logo
  CLASS BLOCK ;
  FOREIGN avali_logo ;
  ORIGIN 0.000 0.000 ;
  SIZE 450.000 BY 528.300 ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal4 ;
        RECT 169.200 362.700 193.500 363.600 ;
        RECT 160.200 361.800 205.200 362.700 ;
        RECT 153.000 360.900 214.200 361.800 ;
        RECT 148.500 360.000 220.500 360.900 ;
        RECT 144.000 359.100 220.500 360.000 ;
        RECT 139.500 358.200 219.600 359.100 ;
        RECT 135.900 357.300 219.600 358.200 ;
        RECT 133.200 356.400 218.700 357.300 ;
        RECT 129.600 355.500 218.700 356.400 ;
        RECT 126.900 354.600 217.800 355.500 ;
        RECT 124.200 353.700 217.800 354.600 ;
        RECT 121.500 352.800 216.900 353.700 ;
        RECT 118.800 351.900 216.000 352.800 ;
        RECT 117.000 351.000 216.000 351.900 ;
        RECT 114.300 350.100 215.100 351.000 ;
        RECT 112.500 349.200 215.100 350.100 ;
        RECT 109.800 348.300 214.200 349.200 ;
        RECT 108.000 347.400 214.200 348.300 ;
        RECT 106.200 346.500 213.300 347.400 ;
        RECT 104.400 345.600 213.300 346.500 ;
        RECT 102.600 344.700 212.400 345.600 ;
        RECT 100.800 343.800 212.400 344.700 ;
        RECT 99.000 342.900 211.500 343.800 ;
        RECT 97.200 342.000 211.500 342.900 ;
        RECT 95.400 341.100 210.600 342.000 ;
        RECT 93.600 340.200 209.700 341.100 ;
        RECT 91.800 339.300 209.700 340.200 ;
        RECT 90.000 338.400 208.800 339.300 ;
        RECT 89.100 337.500 208.800 338.400 ;
        RECT 87.300 336.600 207.900 337.500 ;
        RECT 86.400 335.700 207.900 336.600 ;
        RECT 84.600 334.800 207.000 335.700 ;
        RECT 82.800 333.900 207.000 334.800 ;
        RECT 81.900 333.000 206.100 333.900 ;
        RECT 80.100 332.100 206.100 333.000 ;
        RECT 79.200 331.200 167.400 332.100 ;
        RECT 198.900 331.200 205.200 332.100 ;
        RECT 77.400 330.300 160.200 331.200 ;
        RECT 76.500 329.400 154.800 330.300 ;
        RECT 75.600 328.500 150.300 329.400 ;
        RECT 73.800 327.600 146.700 328.500 ;
        RECT 72.900 326.700 143.100 327.600 ;
        RECT 72.000 325.800 139.500 326.700 ;
        RECT 70.200 324.900 136.800 325.800 ;
        RECT 69.300 324.000 134.100 324.900 ;
        RECT 68.400 323.100 131.400 324.000 ;
        RECT 66.600 322.200 128.700 323.100 ;
        RECT 65.700 321.300 126.900 322.200 ;
        RECT 64.800 320.400 124.200 321.300 ;
        RECT 63.900 319.500 122.400 320.400 ;
        RECT 63.000 318.600 120.600 319.500 ;
        RECT 62.100 317.700 117.900 318.600 ;
        RECT 60.300 316.800 116.100 317.700 ;
        RECT 59.400 315.900 114.300 316.800 ;
        RECT 58.500 315.000 112.500 315.900 ;
        RECT 57.600 314.100 110.700 315.000 ;
        RECT 56.700 313.200 109.800 314.100 ;
        RECT 55.800 312.300 108.000 313.200 ;
        RECT 54.900 311.400 106.200 312.300 ;
        RECT 54.000 310.500 104.400 311.400 ;
        RECT 53.100 309.600 103.500 310.500 ;
        RECT 52.200 308.700 101.700 309.600 ;
        RECT 51.300 307.800 100.800 308.700 ;
        RECT 50.400 306.900 99.000 307.800 ;
        RECT 49.500 306.000 97.200 306.900 ;
        RECT 48.600 305.100 96.300 306.000 ;
        RECT 47.700 304.200 95.400 305.100 ;
        RECT 46.800 303.300 93.600 304.200 ;
        RECT 46.800 302.400 92.700 303.300 ;
        RECT 45.900 301.500 90.900 302.400 ;
        RECT 45.000 300.600 90.000 301.500 ;
        RECT 44.100 299.700 89.100 300.600 ;
        RECT 43.200 298.800 88.200 299.700 ;
        RECT 42.300 297.900 86.400 298.800 ;
        RECT 41.400 297.000 85.500 297.900 ;
        RECT 41.400 296.100 84.600 297.000 ;
        RECT 40.500 295.200 83.700 296.100 ;
        RECT 39.600 294.300 82.800 295.200 ;
        RECT 38.700 293.400 81.900 294.300 ;
        RECT 37.800 292.500 80.100 293.400 ;
        RECT 37.800 291.600 79.200 292.500 ;
        RECT 36.900 290.700 78.300 291.600 ;
        RECT 36.000 289.800 77.400 290.700 ;
        RECT 35.100 288.900 76.500 289.800 ;
        RECT 35.100 288.000 75.600 288.900 ;
        RECT 34.200 287.100 74.700 288.000 ;
        RECT 33.300 286.200 73.800 287.100 ;
        RECT 33.300 285.300 72.900 286.200 ;
        RECT 32.400 284.400 72.000 285.300 ;
        RECT 31.500 283.500 71.100 284.400 ;
        RECT 30.600 281.700 70.200 283.500 ;
        RECT 29.700 280.800 69.300 281.700 ;
        RECT 29.700 279.900 68.400 280.800 ;
        RECT 28.800 279.000 67.500 279.900 ;
        RECT 27.900 278.100 66.600 279.000 ;
        RECT 27.900 277.200 65.700 278.100 ;
        RECT 27.000 276.300 64.800 277.200 ;
        RECT 26.100 275.400 64.800 276.300 ;
        RECT 26.100 274.500 63.900 275.400 ;
        RECT 25.200 273.600 63.000 274.500 ;
        RECT 25.200 272.700 62.100 273.600 ;
        RECT 24.300 271.800 62.100 272.700 ;
        RECT 23.400 270.900 61.200 271.800 ;
        RECT 23.400 270.000 60.300 270.900 ;
        RECT 22.500 268.200 59.400 270.000 ;
        RECT 21.600 267.300 58.500 268.200 ;
        RECT 21.600 266.400 57.600 267.300 ;
        RECT 20.700 265.500 57.600 266.400 ;
        RECT 20.700 264.600 56.700 265.500 ;
        RECT 19.800 262.800 55.800 264.600 ;
        RECT 18.900 261.900 54.900 262.800 ;
        RECT 18.900 261.000 54.000 261.900 ;
        RECT 18.000 260.100 54.000 261.000 ;
        RECT 18.000 259.200 53.100 260.100 ;
        RECT 17.100 257.400 52.200 259.200 ;
        RECT 16.200 255.600 51.300 257.400 ;
        RECT 15.300 253.800 50.400 255.600 ;
        RECT 15.300 252.900 49.500 253.800 ;
        RECT 14.400 252.000 49.500 252.900 ;
        RECT 14.400 251.100 48.600 252.000 ;
        RECT 13.500 250.200 48.600 251.100 ;
        RECT 13.500 249.300 47.700 250.200 ;
        RECT 12.600 248.400 47.700 249.300 ;
        RECT 12.600 246.600 46.800 248.400 ;
        RECT 11.700 244.800 45.900 246.600 ;
        RECT 11.700 243.900 45.000 244.800 ;
        RECT 10.800 243.000 45.000 243.900 ;
        RECT 10.800 242.100 44.100 243.000 ;
        RECT 9.900 241.200 44.100 242.100 ;
        RECT 9.900 239.400 43.200 241.200 ;
        RECT 9.000 236.700 42.300 239.400 ;
        RECT 8.100 234.000 41.400 236.700 ;
        RECT 8.100 233.100 40.500 234.000 ;
        RECT 7.200 232.200 40.500 233.100 ;
        RECT 7.200 230.400 39.600 232.200 ;
        RECT 6.300 229.500 39.600 230.400 ;
        RECT 6.300 226.800 38.700 229.500 ;
        RECT 5.400 223.200 37.800 226.800 ;
        RECT 4.500 220.500 36.900 223.200 ;
        RECT 4.500 218.700 36.000 220.500 ;
        RECT 3.600 216.900 36.000 218.700 ;
        RECT 3.600 214.200 35.100 216.900 ;
        RECT 2.700 212.400 35.100 214.200 ;
        RECT 2.700 208.800 34.200 212.400 ;
        RECT 1.800 207.900 34.200 208.800 ;
        RECT 1.800 202.500 33.300 207.900 ;
        RECT 0.900 201.600 33.300 202.500 ;
        RECT 0.900 193.500 32.400 201.600 ;
        RECT 0.900 191.700 31.500 193.500 ;
        RECT 0.000 171.900 31.500 191.700 ;
        RECT 0.900 170.100 31.500 171.900 ;
        RECT 0.900 161.100 32.400 170.100 ;
        RECT 1.800 155.700 33.300 161.100 ;
        RECT 1.800 154.800 34.200 155.700 ;
        RECT 2.700 151.200 34.200 154.800 ;
        RECT 2.700 149.400 35.100 151.200 ;
        RECT 3.600 146.700 35.100 149.400 ;
        RECT 3.600 144.000 36.000 146.700 ;
        RECT 4.500 143.100 36.000 144.000 ;
        RECT 4.500 140.400 36.900 143.100 ;
        RECT 5.400 136.800 37.800 140.400 ;
        RECT 6.300 134.100 38.700 136.800 ;
        RECT 6.300 133.200 39.600 134.100 ;
        RECT 7.200 131.400 39.600 133.200 ;
        RECT 7.200 130.500 40.500 131.400 ;
        RECT 8.100 129.600 40.500 130.500 ;
        RECT 8.100 126.900 41.400 129.600 ;
        RECT 9.000 124.200 42.300 126.900 ;
        RECT 9.900 122.400 43.200 124.200 ;
        RECT 9.900 121.500 44.100 122.400 ;
        RECT 10.800 120.600 44.100 121.500 ;
        RECT 10.800 119.700 45.000 120.600 ;
        RECT 11.700 118.800 45.000 119.700 ;
        RECT 11.700 117.000 45.900 118.800 ;
        RECT 12.600 116.100 45.900 117.000 ;
        RECT 12.600 114.300 46.800 116.100 ;
        RECT 13.500 112.500 47.700 114.300 ;
        RECT 14.400 110.700 48.600 112.500 ;
        RECT 14.400 109.800 49.500 110.700 ;
        RECT 15.300 108.000 50.400 109.800 ;
        RECT 16.200 106.200 51.300 108.000 ;
        RECT 17.100 104.400 52.200 106.200 ;
        RECT 18.000 103.500 53.100 104.400 ;
        RECT 18.000 102.600 54.000 103.500 ;
        RECT 18.900 101.700 54.000 102.600 ;
        RECT 18.900 100.800 54.900 101.700 ;
        RECT 19.800 99.000 55.800 100.800 ;
        RECT 20.700 97.200 56.700 99.000 ;
        RECT 21.600 96.300 57.600 97.200 ;
        RECT 21.600 95.400 58.500 96.300 ;
        RECT 22.500 93.600 59.400 95.400 ;
        RECT 23.400 92.700 60.300 93.600 ;
        RECT 23.400 91.800 61.200 92.700 ;
        RECT 24.300 90.900 61.200 91.800 ;
        RECT 25.200 90.000 62.100 90.900 ;
        RECT 25.200 89.100 63.000 90.000 ;
        RECT 26.100 88.200 63.900 89.100 ;
        RECT 26.100 87.300 64.800 88.200 ;
        RECT 27.000 86.400 64.800 87.300 ;
        RECT 27.900 85.500 65.700 86.400 ;
        RECT 27.900 84.600 66.600 85.500 ;
        RECT 28.800 83.700 67.500 84.600 ;
        RECT 28.800 82.800 68.400 83.700 ;
        RECT 29.700 81.900 69.300 82.800 ;
        RECT 30.600 81.000 69.300 81.900 ;
        RECT 30.600 80.100 70.200 81.000 ;
        RECT 31.500 79.200 71.100 80.100 ;
        RECT 32.400 78.300 72.000 79.200 ;
        RECT 32.400 77.400 72.900 78.300 ;
        RECT 33.300 76.500 73.800 77.400 ;
        RECT 34.200 75.600 74.700 76.500 ;
        RECT 35.100 74.700 75.600 75.600 ;
        RECT 35.100 73.800 76.500 74.700 ;
        RECT 36.000 72.900 77.400 73.800 ;
        RECT 36.900 72.000 78.300 72.900 ;
        RECT 37.800 71.100 79.200 72.000 ;
        RECT 37.800 70.200 80.100 71.100 ;
        RECT 38.700 69.300 81.000 70.200 ;
        RECT 39.600 68.400 82.800 69.300 ;
        RECT 40.500 67.500 83.700 68.400 ;
        RECT 40.500 66.600 84.600 67.500 ;
        RECT 41.400 65.700 85.500 66.600 ;
        RECT 42.300 64.800 86.400 65.700 ;
        RECT 43.200 63.900 87.300 64.800 ;
        RECT 44.100 63.000 89.100 63.900 ;
        RECT 45.000 62.100 90.000 63.000 ;
        RECT 45.900 61.200 90.900 62.100 ;
        RECT 45.900 60.300 91.800 61.200 ;
        RECT 46.800 59.400 93.600 60.300 ;
        RECT 47.700 58.500 94.500 59.400 ;
        RECT 48.600 57.600 95.400 58.500 ;
        RECT 49.500 56.700 97.200 57.600 ;
        RECT 50.400 55.800 98.100 56.700 ;
        RECT 51.300 54.900 99.900 55.800 ;
        RECT 52.200 54.000 100.800 54.900 ;
        RECT 53.100 53.100 102.600 54.000 ;
        RECT 54.000 52.200 103.500 53.100 ;
        RECT 54.900 51.300 105.300 52.200 ;
        RECT 55.800 50.400 107.100 51.300 ;
        RECT 56.700 49.500 108.900 50.400 ;
        RECT 57.600 48.600 110.700 49.500 ;
        RECT 58.500 47.700 110.700 48.600 ;
        RECT 59.400 46.800 110.700 47.700 ;
        RECT 60.300 45.900 110.700 46.800 ;
        RECT 61.200 45.000 110.700 45.900 ;
        RECT 63.000 44.100 110.700 45.000 ;
        RECT 63.900 43.200 110.700 44.100 ;
        RECT 64.800 42.300 110.700 43.200 ;
        RECT 65.700 41.400 110.700 42.300 ;
        RECT 66.600 40.500 109.800 41.400 ;
        RECT 68.400 39.600 109.800 40.500 ;
        RECT 69.300 38.700 109.800 39.600 ;
        RECT 70.200 37.800 109.800 38.700 ;
        RECT 71.100 36.900 109.800 37.800 ;
        RECT 72.900 36.000 109.800 36.900 ;
        RECT 73.800 35.100 109.800 36.000 ;
        RECT 74.700 34.200 109.800 35.100 ;
        RECT 76.500 33.300 109.800 34.200 ;
        RECT 77.400 32.400 108.900 33.300 ;
        RECT 79.200 31.500 108.900 32.400 ;
        RECT 80.100 30.600 108.900 31.500 ;
        RECT 81.000 29.700 108.900 30.600 ;
        RECT 82.800 28.800 108.900 29.700 ;
        RECT 84.600 27.900 108.900 28.800 ;
        RECT 85.500 27.000 108.900 27.900 ;
        RECT 87.300 26.100 108.900 27.000 ;
        RECT 88.200 25.200 108.000 26.100 ;
        RECT 90.000 24.300 108.000 25.200 ;
        RECT 91.800 23.400 108.000 24.300 ;
        RECT 92.700 22.500 108.000 23.400 ;
        RECT 94.500 21.600 108.000 22.500 ;
        RECT 96.300 20.700 108.000 21.600 ;
        RECT 98.100 19.800 108.000 20.700 ;
        RECT 99.900 18.900 108.000 19.800 ;
        RECT 100.800 18.000 107.100 18.900 ;
        RECT 102.600 17.100 107.100 18.000 ;
        RECT 104.400 16.200 107.100 17.100 ;
        RECT 106.200 15.300 107.100 16.200 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal4 ;
        RECT 352.800 526.500 354.600 527.400 ;
        RECT 351.900 525.600 354.600 526.500 ;
        RECT 351.000 523.800 354.600 525.600 ;
        RECT 350.100 522.900 355.500 523.800 ;
        RECT 349.200 522.000 355.500 522.900 ;
        RECT 348.300 521.100 355.500 522.000 ;
        RECT 347.400 520.200 355.500 521.100 ;
        RECT 346.500 518.400 356.400 520.200 ;
        RECT 345.600 517.500 356.400 518.400 ;
        RECT 344.700 516.600 357.300 517.500 ;
        RECT 343.800 515.700 357.300 516.600 ;
        RECT 342.900 513.900 357.300 515.700 ;
        RECT 342.000 513.000 358.200 513.900 ;
        RECT 341.100 512.100 358.200 513.000 ;
        RECT 340.200 511.200 358.200 512.100 ;
        RECT 339.300 510.300 358.200 511.200 ;
        RECT 338.400 508.500 359.100 510.300 ;
        RECT 337.500 507.600 359.100 508.500 ;
        RECT 336.600 506.700 359.100 507.600 ;
        RECT 335.700 505.800 360.000 506.700 ;
        RECT 334.800 504.000 360.000 505.800 ;
        RECT 333.900 503.100 360.000 504.000 ;
        RECT 333.000 502.200 360.900 503.100 ;
        RECT 332.100 501.300 360.900 502.200 ;
        RECT 331.200 499.500 360.900 501.300 ;
        RECT 330.300 498.600 361.800 499.500 ;
        RECT 329.400 497.700 361.800 498.600 ;
        RECT 328.500 496.800 361.800 497.700 ;
        RECT 327.600 495.900 361.800 496.800 ;
        RECT 327.600 495.000 362.700 495.900 ;
        RECT 326.700 494.100 362.700 495.000 ;
        RECT 325.800 493.200 362.700 494.100 ;
        RECT 324.900 492.300 362.700 493.200 ;
        RECT 324.000 491.400 362.700 492.300 ;
        RECT 324.000 490.500 363.600 491.400 ;
        RECT 323.100 489.600 363.600 490.500 ;
        RECT 322.200 488.700 363.600 489.600 ;
        RECT 321.300 487.800 363.600 488.700 ;
        RECT 320.400 486.900 363.600 487.800 ;
        RECT 320.400 486.000 364.500 486.900 ;
        RECT 319.500 485.100 364.500 486.000 ;
        RECT 318.600 484.200 364.500 485.100 ;
        RECT 317.700 483.300 364.500 484.200 ;
        RECT 316.800 482.400 364.500 483.300 ;
        RECT 316.800 481.500 365.400 482.400 ;
        RECT 315.900 480.600 365.400 481.500 ;
        RECT 315.000 479.700 365.400 480.600 ;
        RECT 314.100 478.800 365.400 479.700 ;
        RECT 313.200 477.000 365.400 478.800 ;
        RECT 312.300 476.100 365.400 477.000 ;
        RECT 311.400 475.200 366.300 476.100 ;
        RECT 310.500 474.300 366.300 475.200 ;
        RECT 309.600 472.500 366.300 474.300 ;
        RECT 308.700 471.600 366.300 472.500 ;
        RECT 307.800 470.700 366.300 471.600 ;
        RECT 306.900 468.900 366.300 470.700 ;
        RECT 306.000 468.000 366.300 468.900 ;
        RECT 305.100 467.100 366.300 468.000 ;
        RECT 304.200 466.200 366.300 467.100 ;
        RECT 303.300 464.400 366.300 466.200 ;
        RECT 302.400 463.500 367.200 464.400 ;
        RECT 301.500 462.600 367.200 463.500 ;
        RECT 300.600 460.800 367.200 462.600 ;
        RECT 299.700 459.900 367.200 460.800 ;
        RECT 298.800 459.000 366.300 459.900 ;
        RECT 297.900 457.200 366.300 459.000 ;
        RECT 297.000 456.300 366.300 457.200 ;
        RECT 296.100 455.400 366.300 456.300 ;
        RECT 295.200 454.500 366.300 455.400 ;
        RECT 294.300 452.700 366.300 454.500 ;
        RECT 293.400 451.800 366.300 452.700 ;
        RECT 292.500 450.900 366.300 451.800 ;
        RECT 291.600 449.100 366.300 450.900 ;
        RECT 290.700 448.200 365.400 449.100 ;
        RECT 289.800 447.300 365.400 448.200 ;
        RECT 288.900 445.500 365.400 447.300 ;
        RECT 288.000 444.600 365.400 445.500 ;
        RECT 287.100 443.700 365.400 444.600 ;
        RECT 286.200 441.900 364.500 443.700 ;
        RECT 285.300 441.000 364.500 441.900 ;
        RECT 284.400 440.100 364.500 441.000 ;
        RECT 283.500 438.300 364.500 440.100 ;
        RECT 282.600 437.400 363.600 438.300 ;
        RECT 281.700 436.500 363.600 437.400 ;
        RECT 280.800 434.700 363.600 436.500 ;
        RECT 279.900 433.800 362.700 434.700 ;
        RECT 279.000 432.000 362.700 433.800 ;
        RECT 278.100 431.100 362.700 432.000 ;
        RECT 277.200 430.200 361.800 431.100 ;
        RECT 276.300 428.400 361.800 430.200 ;
        RECT 275.400 427.500 361.800 428.400 ;
        RECT 274.500 426.600 360.900 427.500 ;
        RECT 273.600 424.800 360.900 426.600 ;
        RECT 272.700 423.900 360.900 424.800 ;
        RECT 271.800 422.100 360.000 423.900 ;
        RECT 270.900 421.200 360.000 422.100 ;
        RECT 270.000 420.300 359.100 421.200 ;
        RECT 269.100 418.500 359.100 420.300 ;
        RECT 268.200 417.600 358.200 418.500 ;
        RECT 267.300 415.800 358.200 417.600 ;
        RECT 266.400 414.900 358.200 415.800 ;
        RECT 265.500 414.000 357.300 414.900 ;
        RECT 264.600 412.200 357.300 414.000 ;
        RECT 263.700 411.300 356.400 412.200 ;
        RECT 262.800 409.500 356.400 411.300 ;
        RECT 261.900 408.600 355.500 409.500 ;
        RECT 261.000 406.800 355.500 408.600 ;
        RECT 260.100 405.900 354.600 406.800 ;
        RECT 259.200 404.100 354.600 405.900 ;
        RECT 258.300 403.200 353.700 404.100 ;
        RECT 257.400 402.300 353.700 403.200 ;
        RECT 256.500 401.400 353.700 402.300 ;
        RECT 256.500 400.500 352.800 401.400 ;
        RECT 255.600 399.600 352.800 400.500 ;
        RECT 254.700 398.700 352.800 399.600 ;
        RECT 254.700 397.800 351.900 398.700 ;
        RECT 253.800 396.900 351.900 397.800 ;
        RECT 252.900 396.000 351.900 396.900 ;
        RECT 252.900 395.100 351.000 396.000 ;
        RECT 252.000 394.200 351.000 395.100 ;
        RECT 251.100 393.300 351.000 394.200 ;
        RECT 251.100 392.400 350.100 393.300 ;
        RECT 250.200 391.500 350.100 392.400 ;
        RECT 249.300 390.600 350.100 391.500 ;
        RECT 249.300 389.700 349.200 390.600 ;
        RECT 248.400 388.800 349.200 389.700 ;
        RECT 247.500 387.000 348.300 388.800 ;
        RECT 246.600 386.100 348.300 387.000 ;
        RECT 245.700 384.300 347.400 386.100 ;
        RECT 244.800 383.400 347.400 384.300 ;
        RECT 244.800 382.500 346.500 383.400 ;
        RECT 243.900 381.600 346.500 382.500 ;
        RECT 243.000 379.800 345.600 381.600 ;
        RECT 242.100 378.900 345.600 379.800 ;
        RECT 241.200 377.100 344.700 378.900 ;
        RECT 240.300 376.200 344.700 377.100 ;
        RECT 239.400 374.400 343.800 376.200 ;
        RECT 238.500 372.600 342.900 374.400 ;
        RECT 237.600 371.700 342.900 372.600 ;
        RECT 236.700 369.900 342.000 371.700 ;
        RECT 235.800 369.000 342.000 369.900 ;
        RECT 234.900 367.200 341.100 369.000 ;
        RECT 234.000 365.400 340.200 367.200 ;
        RECT 233.100 364.500 340.200 365.400 ;
        RECT 232.200 362.700 339.300 364.500 ;
        RECT 231.300 360.900 338.400 362.700 ;
        RECT 230.400 360.000 338.400 360.900 ;
        RECT 229.500 358.200 337.500 360.000 ;
        RECT 228.600 356.400 336.600 358.200 ;
        RECT 227.700 355.500 336.600 356.400 ;
        RECT 226.800 353.700 335.700 355.500 ;
        RECT 225.900 351.900 334.800 353.700 ;
        RECT 225.000 351.000 334.800 351.900 ;
        RECT 224.100 349.200 333.900 351.000 ;
        RECT 223.200 347.400 333.000 349.200 ;
        RECT 222.300 346.500 333.000 347.400 ;
        RECT 222.300 345.600 332.100 346.500 ;
        RECT 221.400 344.700 332.100 345.600 ;
        RECT 221.400 343.800 331.200 344.700 ;
        RECT 220.500 342.900 331.200 343.800 ;
        RECT 219.600 342.000 331.200 342.900 ;
        RECT 219.600 341.100 330.300 342.000 ;
        RECT 218.700 340.200 330.300 341.100 ;
        RECT 218.700 339.300 329.400 340.200 ;
        RECT 217.800 338.400 329.400 339.300 ;
        RECT 217.800 337.500 328.500 338.400 ;
        RECT 216.900 335.700 328.500 337.500 ;
        RECT 216.000 334.800 327.600 335.700 ;
        RECT 215.100 333.900 327.600 334.800 ;
        RECT 215.100 333.000 326.700 333.900 ;
        RECT 214.200 331.200 326.700 333.000 ;
        RECT 213.300 329.400 325.800 331.200 ;
        RECT 212.400 327.600 324.900 329.400 ;
        RECT 211.500 325.800 324.000 327.600 ;
        RECT 210.600 324.900 324.000 325.800 ;
        RECT 210.600 324.000 323.100 324.900 ;
        RECT 209.700 323.100 323.100 324.000 ;
        RECT 209.700 322.200 322.200 323.100 ;
        RECT 208.800 320.400 322.200 322.200 ;
        RECT 207.900 318.600 321.300 320.400 ;
        RECT 207.000 316.800 320.400 318.600 ;
        RECT 206.100 315.000 319.500 316.800 ;
        RECT 205.200 314.100 319.500 315.000 ;
        RECT 205.200 313.200 318.600 314.100 ;
        RECT 204.300 312.300 318.600 313.200 ;
        RECT 204.300 311.400 317.700 312.300 ;
        RECT 203.400 310.500 317.700 311.400 ;
        RECT 203.400 309.600 316.800 310.500 ;
        RECT 202.500 307.800 316.800 309.600 ;
        RECT 201.600 306.000 315.900 307.800 ;
        RECT 200.700 304.200 315.000 306.000 ;
        RECT 199.800 302.400 314.100 304.200 ;
        RECT 198.900 301.500 314.100 302.400 ;
        RECT 198.900 300.600 313.200 301.500 ;
        RECT 198.000 299.700 313.200 300.600 ;
        RECT 198.000 297.900 312.300 299.700 ;
        RECT 197.100 296.100 311.400 297.900 ;
        RECT 196.200 295.200 311.400 296.100 ;
        RECT 196.200 294.300 310.500 295.200 ;
        RECT 195.300 293.400 310.500 294.300 ;
        RECT 195.300 292.500 309.600 293.400 ;
        RECT 194.400 291.600 309.600 292.500 ;
        RECT 194.400 289.800 308.700 291.600 ;
        RECT 193.500 288.900 307.800 289.800 ;
        RECT 193.500 288.000 306.900 288.900 ;
        RECT 192.600 287.100 306.000 288.000 ;
        RECT 192.600 286.200 305.100 287.100 ;
        RECT 191.700 285.300 304.200 286.200 ;
        RECT 191.700 284.400 303.300 285.300 ;
        RECT 190.800 283.500 302.400 284.400 ;
        RECT 190.800 282.600 301.500 283.500 ;
        RECT 190.800 281.700 300.600 282.600 ;
        RECT 189.900 280.800 299.700 281.700 ;
        RECT 189.900 279.900 298.800 280.800 ;
        RECT 189.000 279.000 297.900 279.900 ;
        RECT 189.000 278.100 297.000 279.000 ;
        RECT 189.000 277.200 296.100 278.100 ;
        RECT 188.100 276.300 295.200 277.200 ;
        RECT 188.100 275.400 294.300 276.300 ;
        RECT 187.200 274.500 293.400 275.400 ;
        RECT 187.200 273.600 292.500 274.500 ;
        RECT 186.300 272.700 291.600 273.600 ;
        RECT 186.300 271.800 290.700 272.700 ;
        RECT 186.300 270.900 289.800 271.800 ;
        RECT 185.400 269.100 288.900 270.900 ;
        RECT 184.500 268.200 288.000 269.100 ;
        RECT 184.500 267.300 287.100 268.200 ;
        RECT 184.500 266.400 286.200 267.300 ;
        RECT 183.600 265.500 285.300 266.400 ;
        RECT 183.600 264.600 284.400 265.500 ;
        RECT 182.700 263.700 283.500 264.600 ;
        RECT 182.700 262.800 282.600 263.700 ;
        RECT 182.700 261.900 281.700 262.800 ;
        RECT 181.800 261.000 280.800 261.900 ;
        RECT 181.800 260.100 279.900 261.000 ;
        RECT 180.900 259.200 279.000 260.100 ;
        RECT 180.900 258.300 278.100 259.200 ;
        RECT 180.900 257.400 277.200 258.300 ;
        RECT 180.000 256.500 276.300 257.400 ;
        RECT 180.000 255.600 275.400 256.500 ;
        RECT 179.100 254.700 274.500 255.600 ;
        RECT 179.100 253.800 273.600 254.700 ;
        RECT 179.100 252.900 272.700 253.800 ;
        RECT 178.200 252.000 271.800 252.900 ;
        RECT 178.200 251.100 270.900 252.000 ;
        RECT 178.200 250.200 270.000 251.100 ;
        RECT 177.300 249.300 269.100 250.200 ;
        RECT 177.300 248.400 268.200 249.300 ;
        RECT 176.400 247.500 267.300 248.400 ;
        RECT 176.400 246.600 266.400 247.500 ;
        RECT 176.400 245.700 265.500 246.600 ;
        RECT 175.500 244.800 264.600 245.700 ;
        RECT 175.500 243.900 263.700 244.800 ;
        RECT 175.500 243.000 262.800 243.900 ;
        RECT 174.600 242.100 262.800 243.000 ;
        RECT 174.600 241.200 261.900 242.100 ;
        RECT 173.700 240.300 261.000 241.200 ;
        RECT 173.700 239.400 260.100 240.300 ;
        RECT 173.700 238.500 259.200 239.400 ;
        RECT 172.800 237.600 258.300 238.500 ;
        RECT 172.800 236.700 257.400 237.600 ;
        RECT 172.800 235.800 256.500 236.700 ;
        RECT 171.900 234.900 255.600 235.800 ;
        RECT 171.900 234.000 254.700 234.900 ;
        RECT 171.900 233.100 253.800 234.000 ;
        RECT 171.000 232.200 252.900 233.100 ;
        RECT 171.000 231.300 252.000 232.200 ;
        RECT 170.100 229.500 251.100 231.300 ;
        RECT 170.100 228.600 250.200 229.500 ;
        RECT 169.200 227.700 249.300 228.600 ;
        RECT 169.200 226.800 248.400 227.700 ;
        RECT 169.200 225.900 247.500 226.800 ;
        RECT 168.300 225.000 246.600 225.900 ;
        RECT 168.300 224.100 245.700 225.000 ;
        RECT 168.300 223.200 244.800 224.100 ;
        RECT 167.400 222.300 244.800 223.200 ;
        RECT 167.400 221.400 243.900 222.300 ;
        RECT 167.400 220.500 243.000 221.400 ;
        RECT 166.500 219.600 242.100 220.500 ;
        RECT 166.500 218.700 241.200 219.600 ;
        RECT 166.500 217.800 240.300 218.700 ;
        RECT 165.600 216.000 239.400 217.800 ;
        RECT 165.600 215.100 238.500 216.000 ;
        RECT 164.700 214.200 237.600 215.100 ;
        RECT 164.700 213.300 236.700 214.200 ;
        RECT 164.700 212.400 235.800 213.300 ;
        RECT 163.800 210.600 234.900 212.400 ;
        RECT 163.800 209.700 234.000 210.600 ;
        RECT 162.900 208.800 233.100 209.700 ;
        RECT 162.900 207.900 232.200 208.800 ;
        RECT 162.900 207.000 231.300 207.900 ;
        RECT 162.000 205.200 230.400 207.000 ;
        RECT 162.000 204.300 229.500 205.200 ;
        RECT 161.100 203.400 228.600 204.300 ;
        RECT 161.100 202.500 227.700 203.400 ;
        RECT 161.100 200.700 226.800 202.500 ;
        RECT 160.200 199.800 225.900 200.700 ;
        RECT 160.200 198.900 225.000 199.800 ;
        RECT 160.200 198.000 224.100 198.900 ;
        RECT 159.300 197.100 224.100 198.000 ;
        RECT 159.300 196.200 223.200 197.100 ;
        RECT 159.300 195.300 222.300 196.200 ;
        RECT 158.400 194.400 221.400 195.300 ;
        RECT 158.400 192.600 220.500 194.400 ;
        RECT 157.500 191.700 219.600 192.600 ;
        RECT 157.500 190.800 218.700 191.700 ;
        RECT 157.500 189.900 217.800 190.800 ;
        RECT 156.600 189.000 217.800 189.900 ;
        RECT 156.600 188.100 216.900 189.000 ;
        RECT 156.600 187.200 216.000 188.100 ;
        RECT 156.600 186.300 215.100 187.200 ;
        RECT 155.700 185.400 215.100 186.300 ;
        RECT 155.700 184.500 214.200 185.400 ;
        RECT 155.700 183.600 213.300 184.500 ;
        RECT 154.800 181.800 212.400 183.600 ;
        RECT 154.800 180.900 211.500 181.800 ;
        RECT 153.900 180.000 210.600 180.900 ;
        RECT 153.900 178.200 209.700 180.000 ;
        RECT 153.900 177.300 208.800 178.200 ;
        RECT 153.000 175.500 207.900 177.300 ;
        RECT 153.000 174.600 207.000 175.500 ;
        RECT 152.100 173.700 206.100 174.600 ;
        RECT 152.100 171.900 205.200 173.700 ;
        RECT 152.100 171.000 204.300 171.900 ;
        RECT 151.200 170.100 203.400 171.000 ;
        RECT 151.200 168.300 202.500 170.100 ;
        RECT 150.300 167.400 201.600 168.300 ;
        RECT 150.300 165.600 200.700 167.400 ;
        RECT 149.400 164.700 199.800 165.600 ;
        RECT 149.400 163.800 198.900 164.700 ;
        RECT 149.400 162.000 198.000 163.800 ;
        RECT 148.500 161.100 197.100 162.000 ;
        RECT 148.500 160.200 196.200 161.100 ;
        RECT 148.500 159.300 195.300 160.200 ;
        RECT 147.600 158.400 195.300 159.300 ;
        RECT 147.600 157.500 194.400 158.400 ;
        RECT 147.600 155.700 193.500 157.500 ;
        RECT 146.700 154.800 192.600 155.700 ;
        RECT 146.700 153.000 191.700 154.800 ;
        RECT 145.800 152.100 190.800 153.000 ;
        RECT 145.800 151.200 189.900 152.100 ;
        RECT 145.800 149.400 189.000 151.200 ;
        RECT 144.900 148.500 188.100 149.400 ;
        RECT 144.900 146.700 187.200 148.500 ;
        RECT 144.000 145.800 186.300 146.700 ;
        RECT 144.000 144.000 185.400 145.800 ;
        RECT 144.000 143.100 184.500 144.000 ;
        RECT 143.100 141.300 183.600 143.100 ;
        RECT 143.100 140.400 182.700 141.300 ;
        RECT 142.200 138.600 181.800 140.400 ;
        RECT 142.200 137.700 180.900 138.600 ;
        RECT 142.200 136.800 180.000 137.700 ;
        RECT 141.300 135.900 180.000 136.800 ;
        RECT 141.300 135.000 179.100 135.900 ;
        RECT 141.300 134.100 178.200 135.000 ;
        RECT 140.400 133.200 178.200 134.100 ;
        RECT 140.400 132.300 177.300 133.200 ;
        RECT 140.400 130.500 176.400 132.300 ;
        RECT 139.500 129.600 175.500 130.500 ;
        RECT 139.500 127.800 174.600 129.600 ;
        RECT 138.600 126.900 173.700 127.800 ;
        RECT 138.600 125.100 172.800 126.900 ;
        RECT 138.600 124.200 171.900 125.100 ;
        RECT 137.700 122.400 171.000 124.200 ;
        RECT 137.700 121.500 170.100 122.400 ;
        RECT 137.700 120.600 169.200 121.500 ;
        RECT 136.800 119.700 169.200 120.600 ;
        RECT 136.800 117.900 168.300 119.700 ;
        RECT 136.800 117.000 167.400 117.900 ;
        RECT 135.900 115.200 166.500 117.000 ;
        RECT 135.900 114.300 165.600 115.200 ;
        RECT 135.000 113.400 165.600 114.300 ;
        RECT 135.000 112.500 164.700 113.400 ;
        RECT 135.000 110.700 163.800 112.500 ;
        RECT 134.100 109.800 162.900 110.700 ;
        RECT 134.100 108.000 162.000 109.800 ;
        RECT 134.100 107.100 161.100 108.000 ;
        RECT 133.200 106.200 161.100 107.100 ;
        RECT 133.200 104.400 160.200 106.200 ;
        RECT 133.200 103.500 159.300 104.400 ;
        RECT 132.300 101.700 158.400 103.500 ;
        RECT 132.300 99.900 157.500 101.700 ;
        RECT 131.400 98.100 156.600 99.900 ;
        RECT 131.400 97.200 155.700 98.100 ;
        RECT 131.400 96.300 154.800 97.200 ;
        RECT 130.500 95.400 154.800 96.300 ;
        RECT 130.500 93.600 153.900 95.400 ;
        RECT 130.500 92.700 153.000 93.600 ;
        RECT 129.600 91.800 153.000 92.700 ;
        RECT 129.600 90.000 152.100 91.800 ;
        RECT 129.600 88.200 151.200 90.000 ;
        RECT 128.700 87.300 150.300 88.200 ;
        RECT 128.700 85.500 149.400 87.300 ;
        RECT 128.700 84.600 148.500 85.500 ;
        RECT 127.800 83.700 148.500 84.600 ;
        RECT 127.800 81.900 147.600 83.700 ;
        RECT 127.800 80.100 146.700 81.900 ;
        RECT 126.900 78.300 145.800 80.100 ;
        RECT 126.900 76.500 144.900 78.300 ;
        RECT 126.000 74.700 144.000 76.500 ;
        RECT 126.000 72.900 143.100 74.700 ;
        RECT 126.000 72.000 142.200 72.900 ;
        RECT 125.100 71.100 142.200 72.000 ;
        RECT 125.100 69.300 141.300 71.100 ;
        RECT 125.100 67.500 140.400 69.300 ;
        RECT 124.200 65.700 139.500 67.500 ;
        RECT 124.200 63.900 138.600 65.700 ;
        RECT 124.200 63.000 137.700 63.900 ;
        RECT 123.300 62.100 137.700 63.000 ;
        RECT 123.300 60.300 136.800 62.100 ;
        RECT 123.300 59.400 135.900 60.300 ;
        RECT 122.400 58.500 135.900 59.400 ;
        RECT 122.400 56.700 135.000 58.500 ;
        RECT 122.400 54.900 134.100 56.700 ;
        RECT 121.500 53.100 133.200 54.900 ;
        RECT 121.500 51.300 132.300 53.100 ;
        RECT 121.500 49.500 131.400 51.300 ;
        RECT 120.600 47.700 130.500 49.500 ;
        RECT 120.600 45.900 129.600 47.700 ;
        RECT 120.600 45.000 128.700 45.900 ;
        RECT 119.700 44.100 128.700 45.000 ;
        RECT 119.700 42.300 127.800 44.100 ;
        RECT 119.700 40.500 126.900 42.300 ;
        RECT 118.800 38.700 126.000 40.500 ;
        RECT 118.800 36.900 125.100 38.700 ;
        RECT 118.800 36.000 124.200 36.900 ;
        RECT 117.900 35.100 124.200 36.000 ;
        RECT 117.900 33.300 123.300 35.100 ;
        RECT 117.900 31.500 122.400 33.300 ;
        RECT 117.000 30.600 122.400 31.500 ;
        RECT 117.000 28.800 121.500 30.600 ;
        RECT 117.000 27.000 120.600 28.800 ;
        RECT 117.000 26.100 119.700 27.000 ;
        RECT 116.100 25.200 119.700 26.100 ;
        RECT 116.100 23.400 118.800 25.200 ;
        RECT 116.100 21.600 117.900 23.400 ;
        RECT 115.200 19.800 117.000 21.600 ;
        RECT 115.200 18.000 116.100 19.800 ;
    END
  END vdd
  OBS
      LAYER Metal2 ;
        RECT 0.000 0.000 450.000 528.300 ;
      LAYER Metal3 ;
        RECT 0.000 0.000 450.000 528.300 ;
      LAYER Metal4 ;
        RECT 438.300 376.200 439.200 377.100 ;
        RECT 437.400 375.300 439.200 376.200 ;
        RECT 435.600 374.400 439.200 375.300 ;
        RECT 434.700 373.500 439.200 374.400 ;
        RECT 432.900 372.600 439.200 373.500 ;
        RECT 432.000 371.700 439.200 372.600 ;
        RECT 430.200 370.800 439.200 371.700 ;
        RECT 429.300 369.900 439.200 370.800 ;
        RECT 427.500 369.000 439.200 369.900 ;
        RECT 425.700 368.100 439.200 369.000 ;
        RECT 424.800 367.200 439.200 368.100 ;
        RECT 423.000 366.300 439.200 367.200 ;
        RECT 422.100 365.400 439.200 366.300 ;
        RECT 420.300 364.500 439.200 365.400 ;
        RECT 419.400 363.600 439.200 364.500 ;
        RECT 417.600 362.700 439.200 363.600 ;
        RECT 416.700 361.800 439.200 362.700 ;
        RECT 414.900 360.900 439.200 361.800 ;
        RECT 414.000 360.000 439.200 360.900 ;
        RECT 412.200 359.100 439.200 360.000 ;
        RECT 411.300 358.200 439.200 359.100 ;
        RECT 409.500 357.300 439.200 358.200 ;
        RECT 408.600 356.400 439.200 357.300 ;
        RECT 406.800 355.500 439.200 356.400 ;
        RECT 405.900 354.600 439.200 355.500 ;
        RECT 405.000 353.700 439.200 354.600 ;
        RECT 403.200 352.800 439.200 353.700 ;
        RECT 402.300 351.900 439.200 352.800 ;
        RECT 400.500 351.000 439.200 351.900 ;
        RECT 399.600 350.100 439.200 351.000 ;
        RECT 397.800 349.200 439.200 350.100 ;
        RECT 396.900 348.300 439.200 349.200 ;
        RECT 396.000 347.400 439.200 348.300 ;
        RECT 394.200 346.500 439.200 347.400 ;
        RECT 393.300 345.600 439.200 346.500 ;
        RECT 391.500 344.700 439.200 345.600 ;
        RECT 390.600 343.800 439.200 344.700 ;
        RECT 389.700 342.900 439.200 343.800 ;
        RECT 387.900 342.000 439.200 342.900 ;
        RECT 387.000 341.100 439.200 342.000 ;
        RECT 386.100 340.200 439.200 341.100 ;
        RECT 384.300 339.300 438.300 340.200 ;
        RECT 383.400 338.400 438.300 339.300 ;
        RECT 382.500 337.500 438.300 338.400 ;
        RECT 380.700 336.600 438.300 337.500 ;
        RECT 379.800 335.700 438.300 336.600 ;
        RECT 378.900 334.800 438.300 335.700 ;
        RECT 377.100 333.900 438.300 334.800 ;
        RECT 376.200 333.000 438.300 333.900 ;
        RECT 375.300 332.100 437.400 333.000 ;
        RECT 373.500 331.200 437.400 332.100 ;
        RECT 372.600 330.300 437.400 331.200 ;
        RECT 371.700 329.400 437.400 330.300 ;
        RECT 369.900 328.500 437.400 329.400 ;
        RECT 369.000 327.600 436.500 328.500 ;
        RECT 368.100 326.700 436.500 327.600 ;
        RECT 367.200 325.800 436.500 326.700 ;
        RECT 365.400 324.900 436.500 325.800 ;
        RECT 364.500 324.000 435.600 324.900 ;
        RECT 363.600 323.100 435.600 324.000 ;
        RECT 361.800 322.200 435.600 323.100 ;
        RECT 360.900 321.300 435.600 322.200 ;
        RECT 360.000 320.400 434.700 321.300 ;
        RECT 359.100 319.500 434.700 320.400 ;
        RECT 358.200 318.600 434.700 319.500 ;
        RECT 356.400 317.700 434.700 318.600 ;
        RECT 355.500 316.800 433.800 317.700 ;
        RECT 354.600 315.900 433.800 316.800 ;
        RECT 353.700 315.000 432.900 315.900 ;
        RECT 351.900 314.100 432.900 315.000 ;
        RECT 351.000 313.200 432.000 314.100 ;
        RECT 350.100 312.300 432.000 313.200 ;
        RECT 349.200 311.400 432.000 312.300 ;
        RECT 347.400 310.500 431.100 311.400 ;
        RECT 346.500 309.600 431.100 310.500 ;
        RECT 345.600 308.700 430.200 309.600 ;
        RECT 344.700 307.800 430.200 308.700 ;
        RECT 343.800 306.900 429.300 307.800 ;
        RECT 342.000 306.000 429.300 306.900 ;
        RECT 341.100 305.100 429.300 306.000 ;
        RECT 340.200 304.200 428.400 305.100 ;
        RECT 339.300 303.300 428.400 304.200 ;
        RECT 338.400 302.400 427.500 303.300 ;
        RECT 337.500 301.500 426.600 302.400 ;
        RECT 335.700 300.600 426.600 301.500 ;
        RECT 334.800 299.700 425.700 300.600 ;
        RECT 333.900 298.800 425.700 299.700 ;
        RECT 333.000 297.900 424.800 298.800 ;
        RECT 332.100 297.000 423.900 297.900 ;
        RECT 330.300 296.100 423.900 297.000 ;
        RECT 329.400 295.200 423.000 296.100 ;
        RECT 328.500 294.300 423.000 295.200 ;
        RECT 327.600 293.400 422.100 294.300 ;
        RECT 326.700 292.500 421.200 293.400 ;
        RECT 325.800 291.600 421.200 292.500 ;
        RECT 324.900 290.700 420.300 291.600 ;
        RECT 324.000 289.800 420.300 290.700 ;
        RECT 322.200 288.900 419.400 289.800 ;
        RECT 321.300 288.000 418.500 288.900 ;
        RECT 320.400 287.100 418.500 288.000 ;
        RECT 319.500 286.200 417.600 287.100 ;
        RECT 318.600 285.300 416.700 286.200 ;
        RECT 317.700 284.400 416.700 285.300 ;
        RECT 316.800 283.500 415.800 284.400 ;
        RECT 315.900 282.600 414.900 283.500 ;
        RECT 314.100 281.700 414.000 282.600 ;
        RECT 313.200 280.800 414.000 281.700 ;
        RECT 312.300 279.900 413.100 280.800 ;
        RECT 311.400 279.000 412.200 279.900 ;
        RECT 310.500 278.100 412.200 279.000 ;
        RECT 309.600 277.200 411.300 278.100 ;
        RECT 308.700 276.300 410.400 277.200 ;
        RECT 307.800 275.400 409.500 276.300 ;
        RECT 306.900 274.500 409.500 275.400 ;
        RECT 306.000 273.600 408.600 274.500 ;
        RECT 305.100 272.700 407.700 273.600 ;
        RECT 303.300 271.800 407.700 272.700 ;
        RECT 302.400 270.900 406.800 271.800 ;
        RECT 301.500 270.000 405.900 270.900 ;
        RECT 300.600 269.100 405.000 270.000 ;
        RECT 299.700 268.200 404.100 269.100 ;
        RECT 298.800 267.300 404.100 268.200 ;
        RECT 297.900 266.400 403.200 267.300 ;
        RECT 297.000 265.500 402.300 266.400 ;
        RECT 296.100 264.600 401.400 265.500 ;
        RECT 295.200 263.700 401.400 264.600 ;
        RECT 294.300 262.800 400.500 263.700 ;
        RECT 293.400 261.900 399.600 262.800 ;
        RECT 292.500 261.000 398.700 261.900 ;
        RECT 291.600 260.100 397.800 261.000 ;
        RECT 290.700 259.200 397.800 260.100 ;
        RECT 289.800 258.300 396.900 259.200 ;
        RECT 288.900 257.400 396.000 258.300 ;
        RECT 288.000 256.500 395.100 257.400 ;
        RECT 286.200 255.600 395.100 256.500 ;
        RECT 285.300 254.700 394.200 255.600 ;
        RECT 284.400 253.800 393.300 254.700 ;
        RECT 283.500 252.900 392.400 253.800 ;
        RECT 282.600 252.000 391.500 252.900 ;
        RECT 281.700 251.100 391.500 252.000 ;
        RECT 280.800 250.200 390.600 251.100 ;
        RECT 279.900 249.300 389.700 250.200 ;
        RECT 279.000 248.400 388.800 249.300 ;
        RECT 278.100 247.500 387.900 248.400 ;
        RECT 277.200 246.600 387.900 247.500 ;
        RECT 276.300 245.700 387.000 246.600 ;
        RECT 275.400 244.800 386.100 245.700 ;
        RECT 274.500 243.900 385.200 244.800 ;
        RECT 273.600 243.000 384.300 243.900 ;
        RECT 272.700 242.100 384.300 243.000 ;
        RECT 271.800 241.200 383.400 242.100 ;
        RECT 270.900 240.300 382.500 241.200 ;
        RECT 270.000 239.400 381.600 240.300 ;
        RECT 269.100 238.500 380.700 239.400 ;
        RECT 268.200 237.600 379.800 238.500 ;
        RECT 267.300 236.700 379.800 237.600 ;
        RECT 266.400 235.800 378.900 236.700 ;
        RECT 265.500 234.900 378.000 235.800 ;
        RECT 264.600 234.000 377.100 234.900 ;
        RECT 263.700 233.100 376.200 234.000 ;
        RECT 262.800 232.200 376.200 233.100 ;
        RECT 261.900 231.300 375.300 232.200 ;
        RECT 261.000 230.400 374.400 231.300 ;
        RECT 260.100 229.500 373.500 230.400 ;
        RECT 260.100 228.600 372.600 229.500 ;
        RECT 259.200 227.700 372.600 228.600 ;
        RECT 258.300 226.800 371.700 227.700 ;
        RECT 257.400 225.900 370.800 226.800 ;
        RECT 256.500 225.000 369.900 225.900 ;
        RECT 255.600 224.100 369.000 225.000 ;
        RECT 254.700 223.200 369.000 224.100 ;
        RECT 253.800 222.300 368.100 223.200 ;
        RECT 252.900 221.400 367.200 222.300 ;
        RECT 252.000 220.500 366.300 221.400 ;
        RECT 251.100 219.600 365.400 220.500 ;
        RECT 250.200 218.700 364.500 219.600 ;
        RECT 249.300 217.800 364.500 218.700 ;
        RECT 248.400 216.900 363.600 217.800 ;
        RECT 247.500 216.000 362.700 216.900 ;
        RECT 247.500 215.100 361.800 216.000 ;
        RECT 246.600 214.200 360.900 215.100 ;
        RECT 245.700 213.300 360.900 214.200 ;
        RECT 244.800 212.400 360.000 213.300 ;
        RECT 243.900 211.500 359.100 212.400 ;
        RECT 243.000 210.600 358.200 211.500 ;
        RECT 242.100 209.700 357.300 210.600 ;
        RECT 241.200 208.800 357.300 209.700 ;
        RECT 240.300 207.900 356.400 208.800 ;
        RECT 240.300 207.000 355.500 207.900 ;
        RECT 239.400 206.100 354.600 207.000 ;
        RECT 238.500 205.200 353.700 206.100 ;
        RECT 237.600 204.300 352.800 205.200 ;
        RECT 236.700 203.400 352.800 204.300 ;
        RECT 361.800 203.400 362.700 204.300 ;
        RECT 235.800 202.500 351.900 203.400 ;
        RECT 360.900 202.500 362.700 203.400 ;
        RECT 235.800 201.600 351.000 202.500 ;
        RECT 360.000 201.600 363.600 202.500 ;
        RECT 234.900 200.700 350.100 201.600 ;
        RECT 359.100 200.700 363.600 201.600 ;
        RECT 234.000 199.800 349.200 200.700 ;
        RECT 358.200 199.800 363.600 200.700 ;
        RECT 233.100 198.900 349.200 199.800 ;
        RECT 232.200 198.000 348.300 198.900 ;
        RECT 357.300 198.000 363.600 199.800 ;
        RECT 231.300 197.100 347.400 198.000 ;
        RECT 356.400 197.100 363.600 198.000 ;
        RECT 231.300 196.200 346.500 197.100 ;
        RECT 355.500 196.200 364.500 197.100 ;
        RECT 230.400 195.300 345.600 196.200 ;
        RECT 354.600 195.300 364.500 196.200 ;
        RECT 229.500 194.400 344.700 195.300 ;
        RECT 353.700 194.400 364.500 195.300 ;
        RECT 228.600 193.500 344.700 194.400 ;
        RECT 352.800 193.500 364.500 194.400 ;
        RECT 227.700 192.600 343.800 193.500 ;
        RECT 227.700 191.700 342.900 192.600 ;
        RECT 351.900 191.700 364.500 193.500 ;
        RECT 226.800 190.800 342.000 191.700 ;
        RECT 351.000 190.800 364.500 191.700 ;
        RECT 225.900 189.900 341.100 190.800 ;
        RECT 350.100 189.900 364.500 190.800 ;
        RECT 225.000 189.000 341.100 189.900 ;
        RECT 349.200 189.000 364.500 189.900 ;
        RECT 225.000 188.100 340.200 189.000 ;
        RECT 348.300 188.100 364.500 189.000 ;
        RECT 224.100 187.200 339.300 188.100 ;
        RECT 347.400 187.200 364.500 188.100 ;
        RECT 223.200 186.300 338.400 187.200 ;
        RECT 346.500 186.300 364.500 187.200 ;
        RECT 222.300 185.400 337.500 186.300 ;
        RECT 221.400 184.500 337.500 185.400 ;
        RECT 345.600 184.500 364.500 186.300 ;
        RECT 221.400 183.600 336.600 184.500 ;
        RECT 344.700 183.600 364.500 184.500 ;
        RECT 220.500 182.700 335.700 183.600 ;
        RECT 343.800 182.700 364.500 183.600 ;
        RECT 219.600 181.800 334.800 182.700 ;
        RECT 342.900 181.800 364.500 182.700 ;
        RECT 218.700 180.900 333.900 181.800 ;
        RECT 342.000 180.900 364.500 181.800 ;
        RECT 218.700 180.000 333.000 180.900 ;
        RECT 341.100 180.000 364.500 180.900 ;
        RECT 217.800 179.100 333.000 180.000 ;
        RECT 340.200 179.100 364.500 180.000 ;
        RECT 446.400 179.100 450.000 180.000 ;
        RECT 216.900 178.200 332.100 179.100 ;
        RECT 216.900 177.300 331.200 178.200 ;
        RECT 339.300 177.300 364.500 179.100 ;
        RECT 442.800 178.200 449.100 179.100 ;
        RECT 439.200 177.300 449.100 178.200 ;
        RECT 216.000 176.400 330.300 177.300 ;
        RECT 338.400 176.400 364.500 177.300 ;
        RECT 435.600 176.400 448.200 177.300 ;
        RECT 215.100 175.500 329.400 176.400 ;
        RECT 337.500 175.500 364.500 176.400 ;
        RECT 431.100 175.500 448.200 176.400 ;
        RECT 214.200 174.600 329.400 175.500 ;
        RECT 336.600 174.600 364.500 175.500 ;
        RECT 427.500 174.600 448.200 175.500 ;
        RECT 214.200 173.700 328.500 174.600 ;
        RECT 335.700 173.700 364.500 174.600 ;
        RECT 423.900 173.700 447.300 174.600 ;
        RECT 213.300 172.800 327.600 173.700 ;
        RECT 334.800 172.800 364.500 173.700 ;
        RECT 420.300 172.800 447.300 173.700 ;
        RECT 212.400 171.900 326.700 172.800 ;
        RECT 333.900 171.900 364.500 172.800 ;
        RECT 416.700 171.900 446.400 172.800 ;
        RECT 211.500 171.000 325.800 171.900 ;
        RECT 333.900 171.000 363.600 171.900 ;
        RECT 413.100 171.000 446.400 171.900 ;
        RECT 211.500 170.100 324.900 171.000 ;
        RECT 333.000 170.100 363.600 171.000 ;
        RECT 409.500 170.100 446.400 171.000 ;
        RECT 210.600 169.200 324.900 170.100 ;
        RECT 332.100 169.200 363.600 170.100 ;
        RECT 405.900 169.200 445.500 170.100 ;
        RECT 209.700 168.300 324.000 169.200 ;
        RECT 331.200 168.300 363.600 169.200 ;
        RECT 402.300 168.300 445.500 169.200 ;
        RECT 209.700 167.400 323.100 168.300 ;
        RECT 331.200 167.400 361.800 168.300 ;
        RECT 398.700 167.400 444.600 168.300 ;
        RECT 208.800 166.500 322.200 167.400 ;
        RECT 331.200 166.500 359.100 167.400 ;
        RECT 395.100 166.500 444.600 167.400 ;
        RECT 207.900 164.700 321.300 166.500 ;
        RECT 331.200 165.600 357.300 166.500 ;
        RECT 391.500 165.600 443.700 166.500 ;
        RECT 331.200 164.700 354.600 165.600 ;
        RECT 388.800 164.700 443.700 165.600 ;
        RECT 207.000 163.800 320.400 164.700 ;
        RECT 331.200 163.800 351.900 164.700 ;
        RECT 385.200 163.800 442.800 164.700 ;
        RECT 206.100 162.900 319.500 163.800 ;
        RECT 331.200 162.900 350.100 163.800 ;
        RECT 381.600 162.900 442.800 163.800 ;
        RECT 205.200 162.000 318.600 162.900 ;
        RECT 331.200 162.000 347.400 162.900 ;
        RECT 378.000 162.000 441.900 162.900 ;
        RECT 205.200 161.100 317.700 162.000 ;
        RECT 331.200 161.100 344.700 162.000 ;
        RECT 375.300 161.100 441.900 162.000 ;
        RECT 204.300 160.200 316.800 161.100 ;
        RECT 203.400 159.300 316.800 160.200 ;
        RECT 331.200 160.200 342.000 161.100 ;
        RECT 371.700 160.200 441.000 161.100 ;
        RECT 331.200 159.300 340.200 160.200 ;
        RECT 368.100 159.300 441.000 160.200 ;
        RECT 203.400 158.400 315.900 159.300 ;
        RECT 331.200 158.400 337.500 159.300 ;
        RECT 365.400 158.400 440.100 159.300 ;
        RECT 202.500 157.500 315.000 158.400 ;
        RECT 331.200 157.500 334.800 158.400 ;
        RECT 361.800 157.500 440.100 158.400 ;
        RECT 201.600 156.600 314.100 157.500 ;
        RECT 330.300 156.600 332.100 157.500 ;
        RECT 359.100 156.600 439.200 157.500 ;
        RECT 201.600 155.700 313.200 156.600 ;
        RECT 355.500 155.700 438.300 156.600 ;
        RECT 200.700 154.800 312.300 155.700 ;
        RECT 352.800 154.800 438.300 155.700 ;
        RECT 199.800 153.900 310.500 154.800 ;
        RECT 349.200 153.900 437.400 154.800 ;
        RECT 199.800 153.000 308.700 153.900 ;
        RECT 346.500 153.000 437.400 153.900 ;
        RECT 198.900 152.100 306.900 153.000 ;
        RECT 342.900 152.100 436.500 153.000 ;
        RECT 198.000 151.200 305.100 152.100 ;
        RECT 340.200 151.200 435.600 152.100 ;
        RECT 198.000 150.300 303.300 151.200 ;
        RECT 337.500 150.300 434.700 151.200 ;
        RECT 197.100 149.400 301.500 150.300 ;
        RECT 334.800 149.400 433.800 150.300 ;
        RECT 196.200 148.500 299.700 149.400 ;
        RECT 332.100 148.500 433.800 149.400 ;
        RECT 196.200 147.600 297.900 148.500 ;
        RECT 329.400 147.600 432.900 148.500 ;
        RECT 195.300 146.700 296.100 147.600 ;
        RECT 326.700 146.700 432.000 147.600 ;
        RECT 194.400 145.800 294.300 146.700 ;
        RECT 324.000 145.800 431.100 146.700 ;
        RECT 194.400 144.900 292.500 145.800 ;
        RECT 321.300 144.900 430.200 145.800 ;
        RECT 193.500 144.000 290.700 144.900 ;
        RECT 318.600 144.000 429.300 144.900 ;
        RECT 192.600 143.100 288.900 144.000 ;
        RECT 315.900 143.100 429.300 144.000 ;
        RECT 192.600 142.200 288.000 143.100 ;
        RECT 314.100 142.200 428.400 143.100 ;
        RECT 191.700 141.300 286.200 142.200 ;
        RECT 311.400 141.300 427.500 142.200 ;
        RECT 190.800 140.400 284.400 141.300 ;
        RECT 308.700 140.400 426.600 141.300 ;
        RECT 190.800 139.500 282.600 140.400 ;
        RECT 306.900 139.500 425.700 140.400 ;
        RECT 189.900 138.600 280.800 139.500 ;
        RECT 304.200 138.600 424.800 139.500 ;
        RECT 189.000 137.700 279.000 138.600 ;
        RECT 302.400 137.700 423.900 138.600 ;
        RECT 189.000 136.800 277.200 137.700 ;
        RECT 299.700 136.800 423.000 137.700 ;
        RECT 188.100 135.900 275.400 136.800 ;
        RECT 297.900 135.900 421.200 136.800 ;
        RECT 187.200 135.000 274.500 135.900 ;
        RECT 295.200 135.000 420.300 135.900 ;
        RECT 187.200 134.100 272.700 135.000 ;
        RECT 293.400 134.100 419.400 135.000 ;
        RECT 186.300 133.200 270.900 134.100 ;
        RECT 291.600 133.200 418.500 134.100 ;
        RECT 185.400 132.300 269.100 133.200 ;
        RECT 289.800 132.300 417.600 133.200 ;
        RECT 185.400 131.400 267.300 132.300 ;
        RECT 288.000 131.400 415.800 132.300 ;
        RECT 184.500 130.500 265.500 131.400 ;
        RECT 285.300 130.500 414.900 131.400 ;
        RECT 183.600 129.600 264.600 130.500 ;
        RECT 283.500 129.600 414.000 130.500 ;
        RECT 183.600 128.700 262.800 129.600 ;
        RECT 281.700 128.700 413.100 129.600 ;
        RECT 182.700 127.800 261.000 128.700 ;
        RECT 279.900 127.800 411.300 128.700 ;
        RECT 182.700 126.900 259.200 127.800 ;
        RECT 278.100 126.900 410.400 127.800 ;
        RECT 181.800 126.000 257.400 126.900 ;
        RECT 276.300 126.000 409.500 126.900 ;
        RECT 180.900 125.100 256.500 126.000 ;
        RECT 274.500 125.100 407.700 126.000 ;
        RECT 180.900 124.200 254.700 125.100 ;
        RECT 272.700 124.200 406.800 125.100 ;
        RECT 180.000 123.300 252.900 124.200 ;
        RECT 270.900 123.300 405.000 124.200 ;
        RECT 179.100 122.400 251.100 123.300 ;
        RECT 270.000 122.400 404.100 123.300 ;
        RECT 179.100 121.500 250.200 122.400 ;
        RECT 268.200 121.500 403.200 122.400 ;
        RECT 178.200 120.600 248.400 121.500 ;
        RECT 266.400 120.600 401.400 121.500 ;
        RECT 177.300 119.700 246.600 120.600 ;
        RECT 264.600 119.700 400.500 120.600 ;
        RECT 177.300 118.800 245.700 119.700 ;
        RECT 263.700 118.800 398.700 119.700 ;
        RECT 176.400 117.900 243.900 118.800 ;
        RECT 261.900 117.900 397.800 118.800 ;
        RECT 176.400 117.000 242.100 117.900 ;
        RECT 260.100 117.000 396.000 117.900 ;
        RECT 175.500 116.100 241.200 117.000 ;
        RECT 258.300 116.100 395.100 117.000 ;
        RECT 174.600 115.200 239.400 116.100 ;
        RECT 257.400 115.200 393.300 116.100 ;
        RECT 174.600 114.300 237.600 115.200 ;
        RECT 255.600 114.300 391.500 115.200 ;
        RECT 173.700 113.400 236.700 114.300 ;
        RECT 254.700 113.400 390.600 114.300 ;
        RECT 172.800 112.500 234.900 113.400 ;
        RECT 252.900 112.500 388.800 113.400 ;
        RECT 172.800 111.600 234.000 112.500 ;
        RECT 251.100 111.600 387.900 112.500 ;
        RECT 171.900 110.700 232.200 111.600 ;
        RECT 250.200 110.700 386.100 111.600 ;
        RECT 171.900 109.800 230.400 110.700 ;
        RECT 248.400 109.800 385.200 110.700 ;
        RECT 171.000 108.900 229.500 109.800 ;
        RECT 247.500 108.900 383.400 109.800 ;
        RECT 170.100 108.000 227.700 108.900 ;
        RECT 245.700 108.000 382.500 108.900 ;
        RECT 170.100 107.100 226.800 108.000 ;
        RECT 243.900 107.100 380.700 108.000 ;
        RECT 169.200 106.200 225.000 107.100 ;
        RECT 243.000 106.200 378.900 107.100 ;
        RECT 169.200 105.300 223.200 106.200 ;
        RECT 241.200 105.300 378.000 106.200 ;
        RECT 168.300 104.400 222.300 105.300 ;
        RECT 240.300 104.400 376.200 105.300 ;
        RECT 167.400 103.500 220.500 104.400 ;
        RECT 238.500 103.500 374.400 104.400 ;
        RECT 167.400 102.600 219.600 103.500 ;
        RECT 237.600 102.600 373.500 103.500 ;
        RECT 166.500 101.700 217.800 102.600 ;
        RECT 235.800 101.700 371.700 102.600 ;
        RECT 165.600 100.800 216.900 101.700 ;
        RECT 234.900 100.800 369.900 101.700 ;
        RECT 165.600 99.900 215.100 100.800 ;
        RECT 233.100 99.900 369.000 100.800 ;
        RECT 164.700 99.000 214.200 99.900 ;
        RECT 232.200 99.000 367.200 99.900 ;
        RECT 164.700 98.100 212.400 99.000 ;
        RECT 230.400 98.100 365.400 99.000 ;
        RECT 163.800 97.200 211.500 98.100 ;
        RECT 229.500 97.200 364.500 98.100 ;
        RECT 162.900 96.300 209.700 97.200 ;
        RECT 227.700 96.300 362.700 97.200 ;
        RECT 162.900 95.400 208.800 96.300 ;
        RECT 226.800 95.400 360.900 96.300 ;
        RECT 162.000 94.500 207.000 95.400 ;
        RECT 225.000 94.500 360.000 95.400 ;
        RECT 162.000 93.600 206.100 94.500 ;
        RECT 224.100 93.600 358.200 94.500 ;
        RECT 161.100 92.700 205.200 93.600 ;
        RECT 222.300 92.700 356.400 93.600 ;
        RECT 161.100 91.800 203.400 92.700 ;
        RECT 221.400 91.800 355.500 92.700 ;
        RECT 160.200 90.900 202.500 91.800 ;
        RECT 219.600 90.900 353.700 91.800 ;
        RECT 159.300 90.000 200.700 90.900 ;
        RECT 218.700 90.000 351.900 90.900 ;
        RECT 159.300 89.100 199.800 90.000 ;
        RECT 216.900 89.100 351.000 90.000 ;
        RECT 158.400 88.200 198.000 89.100 ;
        RECT 216.000 88.200 349.200 89.100 ;
        RECT 158.400 87.300 197.100 88.200 ;
        RECT 214.200 87.300 347.400 88.200 ;
        RECT 157.500 86.400 196.200 87.300 ;
        RECT 213.300 86.400 346.500 87.300 ;
        RECT 156.600 85.500 194.400 86.400 ;
        RECT 211.500 85.500 344.700 86.400 ;
        RECT 156.600 84.600 193.500 85.500 ;
        RECT 210.600 84.600 342.900 85.500 ;
        RECT 155.700 83.700 191.700 84.600 ;
        RECT 208.800 83.700 342.000 84.600 ;
        RECT 155.700 82.800 190.800 83.700 ;
        RECT 207.900 82.800 340.200 83.700 ;
        RECT 154.800 81.900 189.900 82.800 ;
        RECT 206.100 81.900 338.400 82.800 ;
        RECT 154.800 81.000 188.100 81.900 ;
        RECT 205.200 81.000 337.500 81.900 ;
        RECT 153.900 80.100 187.200 81.000 ;
        RECT 203.400 80.100 335.700 81.000 ;
        RECT 153.900 79.200 186.300 80.100 ;
        RECT 202.500 79.200 333.900 80.100 ;
        RECT 153.000 78.300 184.500 79.200 ;
        RECT 200.700 78.300 333.000 79.200 ;
        RECT 153.000 77.400 183.600 78.300 ;
        RECT 199.800 77.400 331.200 78.300 ;
        RECT 152.100 76.500 182.700 77.400 ;
        RECT 198.000 76.500 329.400 77.400 ;
        RECT 151.200 75.600 180.900 76.500 ;
        RECT 197.100 75.600 328.500 76.500 ;
        RECT 151.200 74.700 180.000 75.600 ;
        RECT 195.300 74.700 326.700 75.600 ;
        RECT 150.300 73.800 179.100 74.700 ;
        RECT 194.400 73.800 324.900 74.700 ;
        RECT 150.300 72.900 178.200 73.800 ;
        RECT 192.600 72.900 324.000 73.800 ;
        RECT 149.400 72.000 176.400 72.900 ;
        RECT 191.700 72.000 322.200 72.900 ;
        RECT 149.400 71.100 175.500 72.000 ;
        RECT 189.900 71.100 321.300 72.000 ;
        RECT 148.500 70.200 174.600 71.100 ;
        RECT 189.000 70.200 319.500 71.100 ;
        RECT 148.500 69.300 172.800 70.200 ;
        RECT 188.100 69.300 317.700 70.200 ;
        RECT 147.600 68.400 171.900 69.300 ;
        RECT 186.300 68.400 315.900 69.300 ;
        RECT 147.600 67.500 171.000 68.400 ;
        RECT 185.400 67.500 314.100 68.400 ;
        RECT 146.700 66.600 170.100 67.500 ;
        RECT 183.600 66.600 311.400 67.500 ;
        RECT 146.700 65.700 168.300 66.600 ;
        RECT 182.700 65.700 309.600 66.600 ;
        RECT 145.800 64.800 167.400 65.700 ;
        RECT 180.900 64.800 306.900 65.700 ;
        RECT 145.800 63.900 166.500 64.800 ;
        RECT 180.000 63.900 305.100 64.800 ;
        RECT 145.800 63.000 165.600 63.900 ;
        RECT 179.100 63.000 302.400 63.900 ;
        RECT 144.900 62.100 163.800 63.000 ;
        RECT 177.300 62.100 299.700 63.000 ;
        RECT 144.900 61.200 162.900 62.100 ;
        RECT 176.400 61.200 297.900 62.100 ;
        RECT 144.000 60.300 162.000 61.200 ;
        RECT 174.600 60.300 295.200 61.200 ;
        RECT 315.000 60.300 316.800 61.200 ;
        RECT 144.000 59.400 161.100 60.300 ;
        RECT 173.700 59.400 293.400 60.300 ;
        RECT 312.300 59.400 315.900 60.300 ;
        RECT 143.100 58.500 159.300 59.400 ;
        RECT 171.900 58.500 290.700 59.400 ;
        RECT 310.500 58.500 315.000 59.400 ;
        RECT 143.100 57.600 158.400 58.500 ;
        RECT 171.000 57.600 288.900 58.500 ;
        RECT 307.800 57.600 314.100 58.500 ;
        RECT 143.100 56.700 157.500 57.600 ;
        RECT 170.100 56.700 286.200 57.600 ;
        RECT 305.100 56.700 313.200 57.600 ;
        RECT 142.200 55.800 155.700 56.700 ;
        RECT 168.300 55.800 284.400 56.700 ;
        RECT 303.300 55.800 312.300 56.700 ;
        RECT 142.200 54.900 154.800 55.800 ;
        RECT 167.400 54.900 281.700 55.800 ;
        RECT 300.600 54.900 311.400 55.800 ;
        RECT 141.300 54.000 153.900 54.900 ;
        RECT 166.500 54.000 279.900 54.900 ;
        RECT 297.900 54.000 310.500 54.900 ;
        RECT 141.300 53.100 153.000 54.000 ;
        RECT 164.700 53.100 277.200 54.000 ;
        RECT 296.100 53.100 309.600 54.000 ;
        RECT 141.300 52.200 151.200 53.100 ;
        RECT 163.800 52.200 275.400 53.100 ;
        RECT 293.400 52.200 307.800 53.100 ;
        RECT 140.400 51.300 150.300 52.200 ;
        RECT 162.000 51.300 272.700 52.200 ;
        RECT 290.700 51.300 306.900 52.200 ;
        RECT 140.400 50.400 149.400 51.300 ;
        RECT 161.100 50.400 270.000 51.300 ;
        RECT 288.000 50.400 306.000 51.300 ;
        RECT 139.500 49.500 147.600 50.400 ;
        RECT 160.200 49.500 268.200 50.400 ;
        RECT 286.200 49.500 305.100 50.400 ;
        RECT 139.500 48.600 146.700 49.500 ;
        RECT 158.400 48.600 265.500 49.500 ;
        RECT 283.500 48.600 304.200 49.500 ;
        RECT 139.500 47.700 145.800 48.600 ;
        RECT 157.500 47.700 263.700 48.600 ;
        RECT 280.800 47.700 303.300 48.600 ;
        RECT 138.600 46.800 144.000 47.700 ;
        RECT 156.600 46.800 261.000 47.700 ;
        RECT 279.000 46.800 302.400 47.700 ;
        RECT 138.600 45.900 143.100 46.800 ;
        RECT 154.800 45.900 259.200 46.800 ;
        RECT 276.300 45.900 301.500 46.800 ;
        RECT 138.600 45.000 142.200 45.900 ;
        RECT 153.900 45.000 256.500 45.900 ;
        RECT 273.600 45.000 300.600 45.900 ;
        RECT 137.700 44.100 140.400 45.000 ;
        RECT 153.000 44.100 254.700 45.000 ;
        RECT 271.800 44.100 299.700 45.000 ;
        RECT 137.700 43.200 139.500 44.100 ;
        RECT 151.200 43.200 252.000 44.100 ;
        RECT 269.100 43.200 297.900 44.100 ;
        RECT 136.800 42.300 138.600 43.200 ;
        RECT 150.300 42.300 186.300 43.200 ;
        RECT 266.400 42.300 297.000 43.200 ;
        RECT 149.400 41.400 180.000 42.300 ;
        RECT 264.600 41.400 296.100 42.300 ;
        RECT 147.600 40.500 176.400 41.400 ;
        RECT 261.900 40.500 295.200 41.400 ;
        RECT 146.700 39.600 172.800 40.500 ;
        RECT 259.200 39.600 294.300 40.500 ;
        RECT 145.800 38.700 171.000 39.600 ;
        RECT 257.400 38.700 293.400 39.600 ;
        RECT 144.900 37.800 168.300 38.700 ;
        RECT 254.700 37.800 292.500 38.700 ;
        RECT 144.000 36.900 166.500 37.800 ;
        RECT 225.900 36.900 290.700 37.800 ;
        RECT 142.200 36.000 164.700 36.900 ;
        RECT 222.300 36.000 289.800 36.900 ;
        RECT 141.300 35.100 162.000 36.000 ;
        RECT 219.600 35.100 288.900 36.000 ;
        RECT 140.400 34.200 161.100 35.100 ;
        RECT 216.000 34.200 287.100 35.100 ;
        RECT 139.500 33.300 159.300 34.200 ;
        RECT 211.500 33.300 286.200 34.200 ;
        RECT 138.600 32.400 157.500 33.300 ;
        RECT 206.100 32.400 285.300 33.300 ;
        RECT 137.700 31.500 155.700 32.400 ;
        RECT 198.900 31.500 284.400 32.400 ;
        RECT 136.800 30.600 154.800 31.500 ;
        RECT 163.800 30.600 175.500 31.500 ;
        RECT 186.300 30.600 282.600 31.500 ;
        RECT 135.900 29.700 153.000 30.600 ;
        RECT 162.900 29.700 281.700 30.600 ;
        RECT 135.000 28.800 152.100 29.700 ;
        RECT 162.000 28.800 279.900 29.700 ;
        RECT 134.100 27.900 150.300 28.800 ;
        RECT 160.200 27.900 279.000 28.800 ;
        RECT 133.200 27.000 149.400 27.900 ;
        RECT 159.300 27.000 277.200 27.900 ;
        RECT 132.300 26.100 147.600 27.000 ;
        RECT 158.400 26.100 276.300 27.000 ;
        RECT 132.300 25.200 146.700 26.100 ;
        RECT 157.500 25.200 274.500 26.100 ;
        RECT 131.400 24.300 145.800 25.200 ;
        RECT 156.600 24.300 273.600 25.200 ;
        RECT 130.500 23.400 144.000 24.300 ;
        RECT 154.800 23.400 271.800 24.300 ;
        RECT 130.500 22.500 143.100 23.400 ;
        RECT 153.900 22.500 270.000 23.400 ;
        RECT 129.600 21.600 142.200 22.500 ;
        RECT 153.000 21.600 269.100 22.500 ;
        RECT 128.700 20.700 140.400 21.600 ;
        RECT 152.100 20.700 267.300 21.600 ;
        RECT 128.700 19.800 139.500 20.700 ;
        RECT 150.300 19.800 265.500 20.700 ;
        RECT 127.800 18.900 138.600 19.800 ;
        RECT 149.400 18.900 263.700 19.800 ;
        RECT 127.800 18.000 136.800 18.900 ;
        RECT 148.500 18.000 261.900 18.900 ;
        RECT 126.900 17.100 135.900 18.000 ;
        RECT 147.600 17.100 260.100 18.000 ;
        RECT 126.900 16.200 134.100 17.100 ;
        RECT 145.800 16.200 258.300 17.100 ;
        RECT 126.000 15.300 133.200 16.200 ;
        RECT 144.900 15.300 256.500 16.200 ;
        RECT 126.000 14.400 131.400 15.300 ;
        RECT 144.000 14.400 254.700 15.300 ;
        RECT 125.100 13.500 130.500 14.400 ;
        RECT 143.100 13.500 252.000 14.400 ;
        RECT 125.100 12.600 128.700 13.500 ;
        RECT 142.200 12.600 250.200 13.500 ;
        RECT 124.200 11.700 126.900 12.600 ;
        RECT 140.400 11.700 247.500 12.600 ;
        RECT 124.200 10.800 126.000 11.700 ;
        RECT 139.500 10.800 245.700 11.700 ;
        RECT 138.600 9.900 243.000 10.800 ;
        RECT 137.700 9.000 240.300 9.900 ;
        RECT 135.900 8.100 237.600 9.000 ;
        RECT 135.000 7.200 234.900 8.100 ;
        RECT 134.100 6.300 231.300 7.200 ;
        RECT 137.700 5.400 228.600 6.300 ;
        RECT 143.100 4.500 225.000 5.400 ;
        RECT 149.400 3.600 220.500 4.500 ;
        RECT 154.800 2.700 216.900 3.600 ;
        RECT 162.000 1.800 211.500 2.700 ;
        RECT 169.200 0.900 205.200 1.800 ;
        RECT 181.800 0.000 192.600 0.900 ;
  END
END avali_logo
END LIBRARY

