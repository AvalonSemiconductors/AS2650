VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO avali_logo
  CLASS BLOCK ;
  FOREIGN avali_logo ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 352.200 ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal4 ;
        RECT 112.800 241.800 129.000 242.400 ;
        RECT 106.800 241.200 136.800 241.800 ;
        RECT 102.000 240.600 142.800 241.200 ;
        RECT 99.000 240.000 147.000 240.600 ;
        RECT 96.000 239.400 147.000 240.000 ;
        RECT 93.000 238.800 146.400 239.400 ;
        RECT 90.600 238.200 146.400 238.800 ;
        RECT 88.800 237.600 145.800 238.200 ;
        RECT 86.400 237.000 145.800 237.600 ;
        RECT 84.600 236.400 145.200 237.000 ;
        RECT 82.800 235.800 145.200 236.400 ;
        RECT 81.000 235.200 144.600 235.800 ;
        RECT 79.200 234.600 144.000 235.200 ;
        RECT 78.000 234.000 144.000 234.600 ;
        RECT 76.200 233.400 143.400 234.000 ;
        RECT 75.000 232.800 143.400 233.400 ;
        RECT 73.200 232.200 142.800 232.800 ;
        RECT 72.000 231.600 142.800 232.200 ;
        RECT 70.800 231.000 142.200 231.600 ;
        RECT 69.600 230.400 142.200 231.000 ;
        RECT 68.400 229.800 141.600 230.400 ;
        RECT 67.200 229.200 141.600 229.800 ;
        RECT 66.000 228.600 141.000 229.200 ;
        RECT 64.800 228.000 141.000 228.600 ;
        RECT 63.600 227.400 140.400 228.000 ;
        RECT 62.400 226.800 139.800 227.400 ;
        RECT 61.200 226.200 139.800 226.800 ;
        RECT 60.000 225.600 139.200 226.200 ;
        RECT 59.400 225.000 139.200 225.600 ;
        RECT 58.200 224.400 138.600 225.000 ;
        RECT 57.600 223.800 138.600 224.400 ;
        RECT 56.400 223.200 138.000 223.800 ;
        RECT 55.200 222.600 138.000 223.200 ;
        RECT 54.600 222.000 137.400 222.600 ;
        RECT 53.400 221.400 137.400 222.000 ;
        RECT 52.800 220.800 111.600 221.400 ;
        RECT 132.600 220.800 136.800 221.400 ;
        RECT 51.600 220.200 106.800 220.800 ;
        RECT 51.000 219.600 103.200 220.200 ;
        RECT 50.400 219.000 100.200 219.600 ;
        RECT 49.200 218.400 97.800 219.000 ;
        RECT 48.600 217.800 95.400 218.400 ;
        RECT 48.000 217.200 93.000 217.800 ;
        RECT 46.800 216.600 91.200 217.200 ;
        RECT 46.200 216.000 89.400 216.600 ;
        RECT 45.600 215.400 87.600 216.000 ;
        RECT 44.400 214.800 85.800 215.400 ;
        RECT 43.800 214.200 84.600 214.800 ;
        RECT 43.200 213.600 82.800 214.200 ;
        RECT 42.600 213.000 81.600 213.600 ;
        RECT 42.000 212.400 80.400 213.000 ;
        RECT 41.400 211.800 78.600 212.400 ;
        RECT 40.200 211.200 77.400 211.800 ;
        RECT 39.600 210.600 76.200 211.200 ;
        RECT 39.000 210.000 75.000 210.600 ;
        RECT 38.400 209.400 73.800 210.000 ;
        RECT 37.800 208.800 73.200 209.400 ;
        RECT 37.200 208.200 72.000 208.800 ;
        RECT 36.600 207.600 70.800 208.200 ;
        RECT 36.000 207.000 69.600 207.600 ;
        RECT 35.400 206.400 69.000 207.000 ;
        RECT 34.800 205.800 67.800 206.400 ;
        RECT 34.200 205.200 67.200 205.800 ;
        RECT 33.600 204.600 66.000 205.200 ;
        RECT 33.000 204.000 64.800 204.600 ;
        RECT 32.400 203.400 64.200 204.000 ;
        RECT 31.800 202.800 63.600 203.400 ;
        RECT 31.200 202.200 62.400 202.800 ;
        RECT 31.200 201.600 61.800 202.200 ;
        RECT 30.600 201.000 60.600 201.600 ;
        RECT 30.000 200.400 60.000 201.000 ;
        RECT 29.400 199.800 59.400 200.400 ;
        RECT 28.800 199.200 58.800 199.800 ;
        RECT 28.200 198.600 57.600 199.200 ;
        RECT 27.600 198.000 57.000 198.600 ;
        RECT 27.600 197.400 56.400 198.000 ;
        RECT 27.000 196.800 55.800 197.400 ;
        RECT 26.400 196.200 55.200 196.800 ;
        RECT 25.800 195.600 54.600 196.200 ;
        RECT 25.200 195.000 53.400 195.600 ;
        RECT 25.200 194.400 52.800 195.000 ;
        RECT 24.600 193.800 52.200 194.400 ;
        RECT 24.000 193.200 51.600 193.800 ;
        RECT 23.400 192.600 51.000 193.200 ;
        RECT 23.400 192.000 50.400 192.600 ;
        RECT 22.800 191.400 49.800 192.000 ;
        RECT 22.200 190.800 49.200 191.400 ;
        RECT 22.200 190.200 48.600 190.800 ;
        RECT 21.600 189.600 48.000 190.200 ;
        RECT 21.000 189.000 47.400 189.600 ;
        RECT 20.400 187.800 46.800 189.000 ;
        RECT 19.800 187.200 46.200 187.800 ;
        RECT 19.800 186.600 45.600 187.200 ;
        RECT 19.200 186.000 45.000 186.600 ;
        RECT 18.600 185.400 44.400 186.000 ;
        RECT 18.600 184.800 43.800 185.400 ;
        RECT 18.000 184.200 43.200 184.800 ;
        RECT 17.400 183.600 43.200 184.200 ;
        RECT 17.400 183.000 42.600 183.600 ;
        RECT 16.800 182.400 42.000 183.000 ;
        RECT 16.800 181.800 41.400 182.400 ;
        RECT 16.200 181.200 41.400 181.800 ;
        RECT 15.600 180.600 40.800 181.200 ;
        RECT 15.600 180.000 40.200 180.600 ;
        RECT 15.000 178.800 39.600 180.000 ;
        RECT 14.400 178.200 39.000 178.800 ;
        RECT 14.400 177.600 38.400 178.200 ;
        RECT 13.800 177.000 38.400 177.600 ;
        RECT 13.800 176.400 37.800 177.000 ;
        RECT 13.200 175.200 37.200 176.400 ;
        RECT 12.600 174.600 36.600 175.200 ;
        RECT 12.600 174.000 36.000 174.600 ;
        RECT 12.000 173.400 36.000 174.000 ;
        RECT 12.000 172.800 35.400 173.400 ;
        RECT 11.400 171.600 34.800 172.800 ;
        RECT 10.800 170.400 34.200 171.600 ;
        RECT 10.200 169.200 33.600 170.400 ;
        RECT 10.200 168.600 33.000 169.200 ;
        RECT 9.600 168.000 33.000 168.600 ;
        RECT 9.600 167.400 32.400 168.000 ;
        RECT 9.000 166.800 32.400 167.400 ;
        RECT 9.000 166.200 31.800 166.800 ;
        RECT 8.400 165.600 31.800 166.200 ;
        RECT 8.400 164.400 31.200 165.600 ;
        RECT 7.800 163.200 30.600 164.400 ;
        RECT 7.800 162.600 30.000 163.200 ;
        RECT 7.200 162.000 30.000 162.600 ;
        RECT 7.200 161.400 29.400 162.000 ;
        RECT 6.600 160.800 29.400 161.400 ;
        RECT 6.600 159.600 28.800 160.800 ;
        RECT 6.000 157.800 28.200 159.600 ;
        RECT 5.400 156.000 27.600 157.800 ;
        RECT 5.400 155.400 27.000 156.000 ;
        RECT 4.800 154.800 27.000 155.400 ;
        RECT 4.800 153.600 26.400 154.800 ;
        RECT 4.200 153.000 26.400 153.600 ;
        RECT 4.200 151.200 25.800 153.000 ;
        RECT 3.600 148.800 25.200 151.200 ;
        RECT 3.000 147.000 24.600 148.800 ;
        RECT 3.000 145.800 24.000 147.000 ;
        RECT 2.400 144.600 24.000 145.800 ;
        RECT 2.400 142.800 23.400 144.600 ;
        RECT 1.800 141.600 23.400 142.800 ;
        RECT 1.800 139.200 22.800 141.600 ;
        RECT 1.200 138.600 22.800 139.200 ;
        RECT 1.200 135.000 22.200 138.600 ;
        RECT 0.600 134.400 22.200 135.000 ;
        RECT 0.600 129.000 21.600 134.400 ;
        RECT 0.600 127.800 21.000 129.000 ;
        RECT 0.000 114.600 21.000 127.800 ;
        RECT 0.600 113.400 21.000 114.600 ;
        RECT 0.600 107.400 21.600 113.400 ;
        RECT 1.200 103.800 22.200 107.400 ;
        RECT 1.200 103.200 22.800 103.800 ;
        RECT 1.800 100.800 22.800 103.200 ;
        RECT 1.800 99.600 23.400 100.800 ;
        RECT 2.400 97.800 23.400 99.600 ;
        RECT 2.400 96.000 24.000 97.800 ;
        RECT 3.000 95.400 24.000 96.000 ;
        RECT 3.000 93.600 24.600 95.400 ;
        RECT 3.600 91.200 25.200 93.600 ;
        RECT 4.200 89.400 25.800 91.200 ;
        RECT 4.200 88.800 26.400 89.400 ;
        RECT 4.800 87.600 26.400 88.800 ;
        RECT 4.800 87.000 27.000 87.600 ;
        RECT 5.400 86.400 27.000 87.000 ;
        RECT 5.400 84.600 27.600 86.400 ;
        RECT 6.000 82.800 28.200 84.600 ;
        RECT 6.600 81.600 28.800 82.800 ;
        RECT 6.600 81.000 29.400 81.600 ;
        RECT 7.200 80.400 29.400 81.000 ;
        RECT 7.200 79.800 30.000 80.400 ;
        RECT 7.800 79.200 30.000 79.800 ;
        RECT 7.800 78.000 30.600 79.200 ;
        RECT 8.400 77.400 30.600 78.000 ;
        RECT 8.400 76.200 31.200 77.400 ;
        RECT 9.000 75.000 31.800 76.200 ;
        RECT 9.600 73.800 32.400 75.000 ;
        RECT 9.600 73.200 33.000 73.800 ;
        RECT 10.200 72.000 33.600 73.200 ;
        RECT 10.800 70.800 34.200 72.000 ;
        RECT 11.400 69.600 34.800 70.800 ;
        RECT 12.000 69.000 35.400 69.600 ;
        RECT 12.000 68.400 36.000 69.000 ;
        RECT 12.600 67.800 36.000 68.400 ;
        RECT 12.600 67.200 36.600 67.800 ;
        RECT 13.200 66.000 37.200 67.200 ;
        RECT 13.800 64.800 37.800 66.000 ;
        RECT 14.400 64.200 38.400 64.800 ;
        RECT 14.400 63.600 39.000 64.200 ;
        RECT 15.000 62.400 39.600 63.600 ;
        RECT 15.600 61.800 40.200 62.400 ;
        RECT 15.600 61.200 40.800 61.800 ;
        RECT 16.200 60.600 40.800 61.200 ;
        RECT 16.800 60.000 41.400 60.600 ;
        RECT 16.800 59.400 42.000 60.000 ;
        RECT 17.400 58.800 42.600 59.400 ;
        RECT 17.400 58.200 43.200 58.800 ;
        RECT 18.000 57.600 43.200 58.200 ;
        RECT 18.600 57.000 43.800 57.600 ;
        RECT 18.600 56.400 44.400 57.000 ;
        RECT 19.200 55.800 45.000 56.400 ;
        RECT 19.200 55.200 45.600 55.800 ;
        RECT 19.800 54.600 46.200 55.200 ;
        RECT 20.400 54.000 46.200 54.600 ;
        RECT 20.400 53.400 46.800 54.000 ;
        RECT 21.000 52.800 47.400 53.400 ;
        RECT 21.600 52.200 48.000 52.800 ;
        RECT 21.600 51.600 48.600 52.200 ;
        RECT 22.200 51.000 49.200 51.600 ;
        RECT 22.800 50.400 49.800 51.000 ;
        RECT 23.400 49.800 50.400 50.400 ;
        RECT 23.400 49.200 51.000 49.800 ;
        RECT 24.000 48.600 51.600 49.200 ;
        RECT 24.600 48.000 52.200 48.600 ;
        RECT 25.200 47.400 52.800 48.000 ;
        RECT 25.200 46.800 53.400 47.400 ;
        RECT 25.800 46.200 54.000 46.800 ;
        RECT 26.400 45.600 55.200 46.200 ;
        RECT 27.000 45.000 55.800 45.600 ;
        RECT 27.000 44.400 56.400 45.000 ;
        RECT 27.600 43.800 57.000 44.400 ;
        RECT 28.200 43.200 57.600 43.800 ;
        RECT 28.800 42.600 58.200 43.200 ;
        RECT 29.400 42.000 59.400 42.600 ;
        RECT 30.000 41.400 60.000 42.000 ;
        RECT 30.600 40.800 60.600 41.400 ;
        RECT 30.600 40.200 61.200 40.800 ;
        RECT 31.200 39.600 62.400 40.200 ;
        RECT 31.800 39.000 63.000 39.600 ;
        RECT 32.400 38.400 63.600 39.000 ;
        RECT 33.000 37.800 64.800 38.400 ;
        RECT 33.600 37.200 65.400 37.800 ;
        RECT 34.200 36.600 66.600 37.200 ;
        RECT 34.800 36.000 67.200 36.600 ;
        RECT 35.400 35.400 68.400 36.000 ;
        RECT 36.000 34.800 69.000 35.400 ;
        RECT 36.600 34.200 70.200 34.800 ;
        RECT 37.200 33.600 71.400 34.200 ;
        RECT 37.800 33.000 72.600 33.600 ;
        RECT 38.400 32.400 73.800 33.000 ;
        RECT 39.000 31.800 73.800 32.400 ;
        RECT 39.600 31.200 73.800 31.800 ;
        RECT 40.200 30.600 73.800 31.200 ;
        RECT 40.800 30.000 73.800 30.600 ;
        RECT 42.000 29.400 73.800 30.000 ;
        RECT 42.600 28.800 73.800 29.400 ;
        RECT 43.200 28.200 73.800 28.800 ;
        RECT 43.800 27.600 73.800 28.200 ;
        RECT 44.400 27.000 73.200 27.600 ;
        RECT 45.600 26.400 73.200 27.000 ;
        RECT 46.200 25.800 73.200 26.400 ;
        RECT 46.800 25.200 73.200 25.800 ;
        RECT 47.400 24.600 73.200 25.200 ;
        RECT 48.600 24.000 73.200 24.600 ;
        RECT 49.200 23.400 73.200 24.000 ;
        RECT 49.800 22.800 73.200 23.400 ;
        RECT 51.000 22.200 73.200 22.800 ;
        RECT 51.600 21.600 72.600 22.200 ;
        RECT 52.800 21.000 72.600 21.600 ;
        RECT 53.400 20.400 72.600 21.000 ;
        RECT 54.000 19.800 72.600 20.400 ;
        RECT 55.200 19.200 72.600 19.800 ;
        RECT 56.400 18.600 72.600 19.200 ;
        RECT 57.000 18.000 72.600 18.600 ;
        RECT 58.200 17.400 72.600 18.000 ;
        RECT 58.800 16.800 72.000 17.400 ;
        RECT 60.000 16.200 72.000 16.800 ;
        RECT 61.200 15.600 72.000 16.200 ;
        RECT 61.800 15.000 72.000 15.600 ;
        RECT 63.000 14.400 72.000 15.000 ;
        RECT 64.200 13.800 72.000 14.400 ;
        RECT 65.400 13.200 72.000 13.800 ;
        RECT 66.600 12.600 72.000 13.200 ;
        RECT 67.200 12.000 71.400 12.600 ;
        RECT 68.400 11.400 71.400 12.000 ;
        RECT 69.600 10.800 71.400 11.400 ;
        RECT 70.800 10.200 71.400 10.800 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal4 ;
        RECT 235.200 351.000 236.400 351.600 ;
        RECT 234.600 350.400 236.400 351.000 ;
        RECT 234.000 349.200 236.400 350.400 ;
        RECT 233.400 348.600 237.000 349.200 ;
        RECT 232.800 348.000 237.000 348.600 ;
        RECT 232.200 347.400 237.000 348.000 ;
        RECT 231.600 346.800 237.000 347.400 ;
        RECT 231.000 345.600 237.600 346.800 ;
        RECT 230.400 345.000 237.600 345.600 ;
        RECT 229.800 344.400 238.200 345.000 ;
        RECT 229.200 343.800 238.200 344.400 ;
        RECT 228.600 342.600 238.200 343.800 ;
        RECT 228.000 342.000 238.800 342.600 ;
        RECT 227.400 341.400 238.800 342.000 ;
        RECT 226.800 340.800 238.800 341.400 ;
        RECT 226.200 340.200 238.800 340.800 ;
        RECT 225.600 339.000 239.400 340.200 ;
        RECT 225.000 338.400 239.400 339.000 ;
        RECT 224.400 337.800 239.400 338.400 ;
        RECT 223.800 337.200 240.000 337.800 ;
        RECT 223.200 336.000 240.000 337.200 ;
        RECT 222.600 335.400 240.000 336.000 ;
        RECT 222.000 334.800 240.600 335.400 ;
        RECT 221.400 334.200 240.600 334.800 ;
        RECT 220.800 333.000 240.600 334.200 ;
        RECT 220.200 332.400 241.200 333.000 ;
        RECT 219.600 331.800 241.200 332.400 ;
        RECT 219.000 331.200 241.200 331.800 ;
        RECT 218.400 330.600 241.200 331.200 ;
        RECT 218.400 330.000 241.800 330.600 ;
        RECT 217.800 329.400 241.800 330.000 ;
        RECT 217.200 328.800 241.800 329.400 ;
        RECT 216.600 328.200 241.800 328.800 ;
        RECT 216.000 327.600 241.800 328.200 ;
        RECT 216.000 327.000 242.400 327.600 ;
        RECT 215.400 326.400 242.400 327.000 ;
        RECT 214.800 325.800 242.400 326.400 ;
        RECT 214.200 325.200 242.400 325.800 ;
        RECT 213.600 324.600 242.400 325.200 ;
        RECT 213.600 324.000 243.000 324.600 ;
        RECT 213.000 323.400 243.000 324.000 ;
        RECT 212.400 322.800 243.000 323.400 ;
        RECT 211.800 322.200 243.000 322.800 ;
        RECT 211.200 321.600 243.000 322.200 ;
        RECT 211.200 321.000 243.600 321.600 ;
        RECT 210.600 320.400 243.600 321.000 ;
        RECT 210.000 319.800 243.600 320.400 ;
        RECT 209.400 319.200 243.600 319.800 ;
        RECT 208.800 318.000 243.600 319.200 ;
        RECT 208.200 317.400 243.600 318.000 ;
        RECT 207.600 316.800 244.200 317.400 ;
        RECT 207.000 316.200 244.200 316.800 ;
        RECT 206.400 315.000 244.200 316.200 ;
        RECT 205.800 314.400 244.200 315.000 ;
        RECT 205.200 313.800 244.200 314.400 ;
        RECT 204.600 312.600 244.200 313.800 ;
        RECT 204.000 312.000 244.200 312.600 ;
        RECT 203.400 311.400 244.200 312.000 ;
        RECT 202.800 310.800 244.200 311.400 ;
        RECT 202.200 309.600 244.200 310.800 ;
        RECT 201.600 309.000 244.800 309.600 ;
        RECT 201.000 308.400 244.800 309.000 ;
        RECT 200.400 307.200 244.800 308.400 ;
        RECT 199.800 306.600 244.800 307.200 ;
        RECT 199.200 306.000 244.200 306.600 ;
        RECT 198.600 304.800 244.200 306.000 ;
        RECT 198.000 304.200 244.200 304.800 ;
        RECT 197.400 303.600 244.200 304.200 ;
        RECT 196.800 303.000 244.200 303.600 ;
        RECT 196.200 301.800 244.200 303.000 ;
        RECT 195.600 301.200 244.200 301.800 ;
        RECT 195.000 300.600 244.200 301.200 ;
        RECT 194.400 299.400 244.200 300.600 ;
        RECT 193.800 298.800 243.600 299.400 ;
        RECT 193.200 298.200 243.600 298.800 ;
        RECT 192.600 297.000 243.600 298.200 ;
        RECT 192.000 296.400 243.600 297.000 ;
        RECT 191.400 295.800 243.600 296.400 ;
        RECT 190.800 294.600 243.000 295.800 ;
        RECT 190.200 294.000 243.000 294.600 ;
        RECT 189.600 293.400 243.000 294.000 ;
        RECT 189.000 292.200 243.000 293.400 ;
        RECT 188.400 291.600 242.400 292.200 ;
        RECT 187.800 291.000 242.400 291.600 ;
        RECT 187.200 289.800 242.400 291.000 ;
        RECT 186.600 289.200 241.800 289.800 ;
        RECT 186.000 288.000 241.800 289.200 ;
        RECT 185.400 287.400 241.800 288.000 ;
        RECT 184.800 286.800 241.200 287.400 ;
        RECT 184.200 285.600 241.200 286.800 ;
        RECT 183.600 285.000 241.200 285.600 ;
        RECT 183.000 284.400 240.600 285.000 ;
        RECT 182.400 283.200 240.600 284.400 ;
        RECT 181.800 282.600 240.600 283.200 ;
        RECT 181.200 281.400 240.000 282.600 ;
        RECT 180.600 280.800 240.000 281.400 ;
        RECT 180.000 280.200 239.400 280.800 ;
        RECT 179.400 279.000 239.400 280.200 ;
        RECT 178.800 278.400 238.800 279.000 ;
        RECT 178.200 277.200 238.800 278.400 ;
        RECT 177.600 276.600 238.800 277.200 ;
        RECT 177.000 276.000 238.200 276.600 ;
        RECT 176.400 274.800 238.200 276.000 ;
        RECT 175.800 274.200 237.600 274.800 ;
        RECT 175.200 273.000 237.600 274.200 ;
        RECT 174.600 272.400 237.000 273.000 ;
        RECT 174.000 271.200 237.000 272.400 ;
        RECT 173.400 270.600 236.400 271.200 ;
        RECT 172.800 269.400 236.400 270.600 ;
        RECT 172.200 268.800 235.800 269.400 ;
        RECT 171.600 268.200 235.800 268.800 ;
        RECT 171.000 267.600 235.800 268.200 ;
        RECT 171.000 267.000 235.200 267.600 ;
        RECT 170.400 266.400 235.200 267.000 ;
        RECT 169.800 265.800 235.200 266.400 ;
        RECT 169.800 265.200 234.600 265.800 ;
        RECT 169.200 264.600 234.600 265.200 ;
        RECT 168.600 264.000 234.600 264.600 ;
        RECT 168.600 263.400 234.000 264.000 ;
        RECT 168.000 262.800 234.000 263.400 ;
        RECT 167.400 262.200 234.000 262.800 ;
        RECT 167.400 261.600 233.400 262.200 ;
        RECT 166.800 261.000 233.400 261.600 ;
        RECT 166.200 260.400 233.400 261.000 ;
        RECT 166.200 259.800 232.800 260.400 ;
        RECT 165.600 259.200 232.800 259.800 ;
        RECT 165.000 258.000 232.200 259.200 ;
        RECT 164.400 257.400 232.200 258.000 ;
        RECT 163.800 256.200 231.600 257.400 ;
        RECT 163.200 255.600 231.600 256.200 ;
        RECT 163.200 255.000 231.000 255.600 ;
        RECT 162.600 254.400 231.000 255.000 ;
        RECT 162.000 253.200 230.400 254.400 ;
        RECT 161.400 252.600 230.400 253.200 ;
        RECT 160.800 251.400 229.800 252.600 ;
        RECT 160.200 250.800 229.800 251.400 ;
        RECT 159.600 249.600 229.200 250.800 ;
        RECT 159.000 248.400 228.600 249.600 ;
        RECT 158.400 247.800 228.600 248.400 ;
        RECT 157.800 246.600 228.000 247.800 ;
        RECT 157.200 246.000 228.000 246.600 ;
        RECT 156.600 244.800 227.400 246.000 ;
        RECT 156.000 243.600 226.800 244.800 ;
        RECT 155.400 243.000 226.800 243.600 ;
        RECT 154.800 241.800 226.200 243.000 ;
        RECT 154.200 240.600 225.600 241.800 ;
        RECT 153.600 240.000 225.600 240.600 ;
        RECT 153.000 238.800 225.000 240.000 ;
        RECT 152.400 237.600 224.400 238.800 ;
        RECT 151.800 237.000 224.400 237.600 ;
        RECT 151.200 235.800 223.800 237.000 ;
        RECT 150.600 234.600 223.200 235.800 ;
        RECT 150.000 234.000 223.200 234.600 ;
        RECT 149.400 232.800 222.600 234.000 ;
        RECT 148.800 231.600 222.000 232.800 ;
        RECT 148.200 231.000 222.000 231.600 ;
        RECT 148.200 230.400 221.400 231.000 ;
        RECT 147.600 229.800 221.400 230.400 ;
        RECT 147.600 229.200 220.800 229.800 ;
        RECT 147.000 228.600 220.800 229.200 ;
        RECT 146.400 228.000 220.800 228.600 ;
        RECT 146.400 227.400 220.200 228.000 ;
        RECT 145.800 226.800 220.200 227.400 ;
        RECT 145.800 226.200 219.600 226.800 ;
        RECT 145.200 225.600 219.600 226.200 ;
        RECT 145.200 225.000 219.000 225.600 ;
        RECT 144.600 223.800 219.000 225.000 ;
        RECT 144.000 223.200 218.400 223.800 ;
        RECT 143.400 222.600 218.400 223.200 ;
        RECT 143.400 222.000 217.800 222.600 ;
        RECT 142.800 220.800 217.800 222.000 ;
        RECT 142.200 219.600 217.200 220.800 ;
        RECT 141.600 218.400 216.600 219.600 ;
        RECT 141.000 217.200 216.000 218.400 ;
        RECT 140.400 216.600 216.000 217.200 ;
        RECT 140.400 216.000 215.400 216.600 ;
        RECT 139.800 215.400 215.400 216.000 ;
        RECT 139.800 214.800 214.800 215.400 ;
        RECT 139.200 213.600 214.800 214.800 ;
        RECT 138.600 212.400 214.200 213.600 ;
        RECT 138.000 211.200 213.600 212.400 ;
        RECT 137.400 210.000 213.000 211.200 ;
        RECT 136.800 209.400 213.000 210.000 ;
        RECT 136.800 208.800 212.400 209.400 ;
        RECT 136.200 208.200 212.400 208.800 ;
        RECT 136.200 207.600 211.800 208.200 ;
        RECT 135.600 207.000 211.800 207.600 ;
        RECT 135.600 206.400 211.200 207.000 ;
        RECT 135.000 205.200 211.200 206.400 ;
        RECT 134.400 204.000 210.600 205.200 ;
        RECT 133.800 202.800 210.000 204.000 ;
        RECT 133.200 201.600 209.400 202.800 ;
        RECT 132.600 201.000 209.400 201.600 ;
        RECT 132.600 200.400 208.800 201.000 ;
        RECT 132.000 199.800 208.800 200.400 ;
        RECT 132.000 198.600 208.200 199.800 ;
        RECT 131.400 197.400 207.600 198.600 ;
        RECT 130.800 196.800 207.600 197.400 ;
        RECT 130.800 196.200 207.000 196.800 ;
        RECT 130.200 195.600 207.000 196.200 ;
        RECT 130.200 195.000 206.400 195.600 ;
        RECT 129.600 194.400 206.400 195.000 ;
        RECT 129.600 193.200 205.800 194.400 ;
        RECT 129.000 192.600 205.200 193.200 ;
        RECT 129.000 192.000 204.600 192.600 ;
        RECT 128.400 191.400 204.000 192.000 ;
        RECT 128.400 190.800 203.400 191.400 ;
        RECT 127.800 190.200 202.800 190.800 ;
        RECT 127.800 189.600 202.200 190.200 ;
        RECT 127.200 189.000 201.600 189.600 ;
        RECT 127.200 188.400 201.000 189.000 ;
        RECT 127.200 187.800 200.400 188.400 ;
        RECT 126.600 187.200 199.800 187.800 ;
        RECT 126.600 186.600 199.200 187.200 ;
        RECT 126.000 186.000 198.600 186.600 ;
        RECT 126.000 185.400 198.000 186.000 ;
        RECT 126.000 184.800 197.400 185.400 ;
        RECT 125.400 184.200 196.800 184.800 ;
        RECT 125.400 183.600 196.200 184.200 ;
        RECT 124.800 183.000 195.600 183.600 ;
        RECT 124.800 182.400 195.000 183.000 ;
        RECT 124.200 181.800 194.400 182.400 ;
        RECT 124.200 181.200 193.800 181.800 ;
        RECT 124.200 180.600 193.200 181.200 ;
        RECT 123.600 179.400 192.600 180.600 ;
        RECT 123.000 178.800 192.000 179.400 ;
        RECT 123.000 178.200 191.400 178.800 ;
        RECT 123.000 177.600 190.800 178.200 ;
        RECT 122.400 177.000 190.200 177.600 ;
        RECT 122.400 176.400 189.600 177.000 ;
        RECT 121.800 175.800 189.000 176.400 ;
        RECT 121.800 175.200 188.400 175.800 ;
        RECT 121.800 174.600 187.800 175.200 ;
        RECT 121.200 174.000 187.200 174.600 ;
        RECT 121.200 173.400 186.600 174.000 ;
        RECT 120.600 172.800 186.000 173.400 ;
        RECT 120.600 172.200 185.400 172.800 ;
        RECT 120.600 171.600 184.800 172.200 ;
        RECT 120.000 171.000 184.200 171.600 ;
        RECT 120.000 170.400 183.600 171.000 ;
        RECT 119.400 169.800 183.000 170.400 ;
        RECT 119.400 169.200 182.400 169.800 ;
        RECT 119.400 168.600 181.800 169.200 ;
        RECT 118.800 168.000 181.200 168.600 ;
        RECT 118.800 167.400 180.600 168.000 ;
        RECT 118.800 166.800 180.000 167.400 ;
        RECT 118.200 166.200 179.400 166.800 ;
        RECT 118.200 165.600 178.800 166.200 ;
        RECT 117.600 165.000 178.200 165.600 ;
        RECT 117.600 164.400 177.600 165.000 ;
        RECT 117.600 163.800 177.000 164.400 ;
        RECT 117.000 163.200 176.400 163.800 ;
        RECT 117.000 162.600 175.800 163.200 ;
        RECT 117.000 162.000 175.200 162.600 ;
        RECT 116.400 161.400 175.200 162.000 ;
        RECT 116.400 160.800 174.600 161.400 ;
        RECT 115.800 160.200 174.000 160.800 ;
        RECT 115.800 159.600 173.400 160.200 ;
        RECT 115.800 159.000 172.800 159.600 ;
        RECT 115.200 158.400 172.200 159.000 ;
        RECT 115.200 157.800 171.600 158.400 ;
        RECT 115.200 157.200 171.000 157.800 ;
        RECT 114.600 156.600 170.400 157.200 ;
        RECT 114.600 156.000 169.800 156.600 ;
        RECT 114.600 155.400 169.200 156.000 ;
        RECT 114.000 154.800 168.600 155.400 ;
        RECT 114.000 154.200 168.000 154.800 ;
        RECT 113.400 153.000 167.400 154.200 ;
        RECT 113.400 152.400 166.800 153.000 ;
        RECT 112.800 151.800 166.200 152.400 ;
        RECT 112.800 151.200 165.600 151.800 ;
        RECT 112.800 150.600 165.000 151.200 ;
        RECT 112.200 150.000 164.400 150.600 ;
        RECT 112.200 149.400 163.800 150.000 ;
        RECT 112.200 148.800 163.200 149.400 ;
        RECT 111.600 148.200 163.200 148.800 ;
        RECT 111.600 147.600 162.600 148.200 ;
        RECT 111.600 147.000 162.000 147.600 ;
        RECT 111.000 146.400 161.400 147.000 ;
        RECT 111.000 145.800 160.800 146.400 ;
        RECT 111.000 145.200 160.200 145.800 ;
        RECT 110.400 144.000 159.600 145.200 ;
        RECT 110.400 143.400 159.000 144.000 ;
        RECT 109.800 142.800 158.400 143.400 ;
        RECT 109.800 142.200 157.800 142.800 ;
        RECT 109.800 141.600 157.200 142.200 ;
        RECT 109.200 140.400 156.600 141.600 ;
        RECT 109.200 139.800 156.000 140.400 ;
        RECT 108.600 139.200 155.400 139.800 ;
        RECT 108.600 138.600 154.800 139.200 ;
        RECT 108.600 138.000 154.200 138.600 ;
        RECT 108.000 136.800 153.600 138.000 ;
        RECT 108.000 136.200 153.000 136.800 ;
        RECT 107.400 135.600 152.400 136.200 ;
        RECT 107.400 135.000 151.800 135.600 ;
        RECT 107.400 133.800 151.200 135.000 ;
        RECT 106.800 133.200 150.600 133.800 ;
        RECT 106.800 132.600 150.000 133.200 ;
        RECT 106.800 132.000 149.400 132.600 ;
        RECT 106.200 131.400 149.400 132.000 ;
        RECT 106.200 130.800 148.800 131.400 ;
        RECT 106.200 130.200 148.200 130.800 ;
        RECT 105.600 129.600 147.600 130.200 ;
        RECT 105.600 128.400 147.000 129.600 ;
        RECT 105.000 127.800 146.400 128.400 ;
        RECT 105.000 127.200 145.800 127.800 ;
        RECT 105.000 126.600 145.200 127.200 ;
        RECT 104.400 126.000 145.200 126.600 ;
        RECT 104.400 125.400 144.600 126.000 ;
        RECT 104.400 124.800 144.000 125.400 ;
        RECT 104.400 124.200 143.400 124.800 ;
        RECT 103.800 123.600 143.400 124.200 ;
        RECT 103.800 123.000 142.800 123.600 ;
        RECT 103.800 122.400 142.200 123.000 ;
        RECT 103.200 121.200 141.600 122.400 ;
        RECT 103.200 120.600 141.000 121.200 ;
        RECT 102.600 120.000 140.400 120.600 ;
        RECT 102.600 118.800 139.800 120.000 ;
        RECT 102.600 118.200 139.200 118.800 ;
        RECT 102.000 117.000 138.600 118.200 ;
        RECT 102.000 116.400 138.000 117.000 ;
        RECT 101.400 115.800 137.400 116.400 ;
        RECT 101.400 114.600 136.800 115.800 ;
        RECT 101.400 114.000 136.200 114.600 ;
        RECT 100.800 113.400 135.600 114.000 ;
        RECT 100.800 112.200 135.000 113.400 ;
        RECT 100.200 111.600 134.400 112.200 ;
        RECT 100.200 110.400 133.800 111.600 ;
        RECT 99.600 109.800 133.200 110.400 ;
        RECT 99.600 109.200 132.600 109.800 ;
        RECT 99.600 108.000 132.000 109.200 ;
        RECT 99.000 107.400 131.400 108.000 ;
        RECT 99.000 106.800 130.800 107.400 ;
        RECT 99.000 106.200 130.200 106.800 ;
        RECT 98.400 105.600 130.200 106.200 ;
        RECT 98.400 105.000 129.600 105.600 ;
        RECT 98.400 103.800 129.000 105.000 ;
        RECT 97.800 103.200 128.400 103.800 ;
        RECT 97.800 102.000 127.800 103.200 ;
        RECT 97.200 101.400 127.200 102.000 ;
        RECT 97.200 100.800 126.600 101.400 ;
        RECT 97.200 99.600 126.000 100.800 ;
        RECT 96.600 99.000 125.400 99.600 ;
        RECT 96.600 97.800 124.800 99.000 ;
        RECT 96.000 97.200 124.200 97.800 ;
        RECT 96.000 96.000 123.600 97.200 ;
        RECT 96.000 95.400 123.000 96.000 ;
        RECT 95.400 94.200 122.400 95.400 ;
        RECT 95.400 93.600 121.800 94.200 ;
        RECT 94.800 92.400 121.200 93.600 ;
        RECT 94.800 91.800 120.600 92.400 ;
        RECT 94.800 91.200 120.000 91.800 ;
        RECT 94.200 90.600 120.000 91.200 ;
        RECT 94.200 90.000 119.400 90.600 ;
        RECT 94.200 89.400 118.800 90.000 ;
        RECT 93.600 88.800 118.800 89.400 ;
        RECT 93.600 88.200 118.200 88.800 ;
        RECT 93.600 87.000 117.600 88.200 ;
        RECT 93.000 86.400 117.000 87.000 ;
        RECT 93.000 85.200 116.400 86.400 ;
        RECT 92.400 84.600 115.800 85.200 ;
        RECT 92.400 83.400 115.200 84.600 ;
        RECT 92.400 82.800 114.600 83.400 ;
        RECT 91.800 81.600 114.000 82.800 ;
        RECT 91.800 81.000 113.400 81.600 ;
        RECT 91.800 80.400 112.800 81.000 ;
        RECT 91.200 79.800 112.800 80.400 ;
        RECT 91.200 78.600 112.200 79.800 ;
        RECT 91.200 78.000 111.600 78.600 ;
        RECT 90.600 76.800 111.000 78.000 ;
        RECT 90.600 76.200 110.400 76.800 ;
        RECT 90.000 75.600 110.400 76.200 ;
        RECT 90.000 75.000 109.800 75.600 ;
        RECT 90.000 73.800 109.200 75.000 ;
        RECT 89.400 73.200 108.600 73.800 ;
        RECT 89.400 72.000 108.000 73.200 ;
        RECT 89.400 71.400 107.400 72.000 ;
        RECT 88.800 70.800 107.400 71.400 ;
        RECT 88.800 69.600 106.800 70.800 ;
        RECT 88.800 69.000 106.200 69.600 ;
        RECT 88.200 67.800 105.600 69.000 ;
        RECT 88.200 66.600 105.000 67.800 ;
        RECT 87.600 65.400 104.400 66.600 ;
        RECT 87.600 64.800 103.800 65.400 ;
        RECT 87.600 64.200 103.200 64.800 ;
        RECT 87.000 63.600 103.200 64.200 ;
        RECT 87.000 62.400 102.600 63.600 ;
        RECT 87.000 61.800 102.000 62.400 ;
        RECT 86.400 61.200 102.000 61.800 ;
        RECT 86.400 60.000 101.400 61.200 ;
        RECT 86.400 58.800 100.800 60.000 ;
        RECT 85.800 58.200 100.200 58.800 ;
        RECT 85.800 57.000 99.600 58.200 ;
        RECT 85.800 56.400 99.000 57.000 ;
        RECT 85.200 55.800 99.000 56.400 ;
        RECT 85.200 54.600 98.400 55.800 ;
        RECT 85.200 53.400 97.800 54.600 ;
        RECT 84.600 52.200 97.200 53.400 ;
        RECT 84.600 51.000 96.600 52.200 ;
        RECT 84.000 49.800 96.000 51.000 ;
        RECT 84.000 48.600 95.400 49.800 ;
        RECT 84.000 48.000 94.800 48.600 ;
        RECT 83.400 47.400 94.800 48.000 ;
        RECT 83.400 46.200 94.200 47.400 ;
        RECT 83.400 45.000 93.600 46.200 ;
        RECT 82.800 43.800 93.000 45.000 ;
        RECT 82.800 42.600 92.400 43.800 ;
        RECT 82.800 42.000 91.800 42.600 ;
        RECT 82.200 41.400 91.800 42.000 ;
        RECT 82.200 40.200 91.200 41.400 ;
        RECT 82.200 39.600 90.600 40.200 ;
        RECT 81.600 39.000 90.600 39.600 ;
        RECT 81.600 37.800 90.000 39.000 ;
        RECT 81.600 36.600 89.400 37.800 ;
        RECT 81.000 35.400 88.800 36.600 ;
        RECT 81.000 34.200 88.200 35.400 ;
        RECT 81.000 33.000 87.600 34.200 ;
        RECT 80.400 31.800 87.000 33.000 ;
        RECT 80.400 30.600 86.400 31.800 ;
        RECT 80.400 30.000 85.800 30.600 ;
        RECT 79.800 29.400 85.800 30.000 ;
        RECT 79.800 28.200 85.200 29.400 ;
        RECT 79.800 27.000 84.600 28.200 ;
        RECT 79.200 25.800 84.000 27.000 ;
        RECT 79.200 24.600 83.400 25.800 ;
        RECT 79.200 24.000 82.800 24.600 ;
        RECT 78.600 23.400 82.800 24.000 ;
        RECT 78.600 22.200 82.200 23.400 ;
        RECT 78.600 21.000 81.600 22.200 ;
        RECT 78.000 20.400 81.600 21.000 ;
        RECT 78.000 19.200 81.000 20.400 ;
        RECT 78.000 18.000 80.400 19.200 ;
        RECT 78.000 17.400 79.800 18.000 ;
        RECT 77.400 16.800 79.800 17.400 ;
        RECT 77.400 15.600 79.200 16.800 ;
        RECT 77.400 14.400 78.600 15.600 ;
        RECT 76.800 13.200 78.000 14.400 ;
        RECT 76.800 12.000 77.400 13.200 ;
    END
  END vdd
  OBS
      LAYER Metal2 ;
        RECT 0.000 0.000 300.000 352.200 ;
      LAYER Metal3 ;
        RECT 0.000 0.000 300.000 352.200 ;
      LAYER Metal4 ;
        RECT 292.200 250.800 292.800 251.400 ;
        RECT 291.600 250.200 292.800 250.800 ;
        RECT 290.400 249.600 292.800 250.200 ;
        RECT 289.800 249.000 292.800 249.600 ;
        RECT 288.600 248.400 292.800 249.000 ;
        RECT 288.000 247.800 292.800 248.400 ;
        RECT 286.800 247.200 292.800 247.800 ;
        RECT 286.200 246.600 292.800 247.200 ;
        RECT 285.000 246.000 292.800 246.600 ;
        RECT 283.800 245.400 292.800 246.000 ;
        RECT 283.200 244.800 292.800 245.400 ;
        RECT 282.000 244.200 292.800 244.800 ;
        RECT 281.400 243.600 292.800 244.200 ;
        RECT 280.200 243.000 292.800 243.600 ;
        RECT 279.600 242.400 292.800 243.000 ;
        RECT 278.400 241.800 292.800 242.400 ;
        RECT 277.800 241.200 292.800 241.800 ;
        RECT 276.600 240.600 292.800 241.200 ;
        RECT 276.000 240.000 292.800 240.600 ;
        RECT 274.800 239.400 292.800 240.000 ;
        RECT 274.200 238.800 292.800 239.400 ;
        RECT 273.000 238.200 292.800 238.800 ;
        RECT 272.400 237.600 292.800 238.200 ;
        RECT 271.200 237.000 292.800 237.600 ;
        RECT 270.600 236.400 292.800 237.000 ;
        RECT 270.000 235.800 292.800 236.400 ;
        RECT 268.800 235.200 292.800 235.800 ;
        RECT 268.200 234.600 292.800 235.200 ;
        RECT 267.000 234.000 292.800 234.600 ;
        RECT 266.400 233.400 292.800 234.000 ;
        RECT 265.200 232.800 292.800 233.400 ;
        RECT 264.600 232.200 292.800 232.800 ;
        RECT 264.000 231.600 292.800 232.200 ;
        RECT 262.800 231.000 292.800 231.600 ;
        RECT 262.200 230.400 292.800 231.000 ;
        RECT 261.000 229.800 292.800 230.400 ;
        RECT 260.400 229.200 292.800 229.800 ;
        RECT 259.800 228.600 292.800 229.200 ;
        RECT 258.600 228.000 292.800 228.600 ;
        RECT 258.000 227.400 292.800 228.000 ;
        RECT 257.400 226.800 292.800 227.400 ;
        RECT 256.200 226.200 292.200 226.800 ;
        RECT 255.600 225.600 292.200 226.200 ;
        RECT 255.000 225.000 292.200 225.600 ;
        RECT 253.800 224.400 292.200 225.000 ;
        RECT 253.200 223.800 292.200 224.400 ;
        RECT 252.600 223.200 292.200 223.800 ;
        RECT 251.400 222.600 292.200 223.200 ;
        RECT 250.800 222.000 292.200 222.600 ;
        RECT 250.200 221.400 291.600 222.000 ;
        RECT 249.000 220.800 291.600 221.400 ;
        RECT 248.400 220.200 291.600 220.800 ;
        RECT 247.800 219.600 291.600 220.200 ;
        RECT 246.600 219.000 291.600 219.600 ;
        RECT 246.000 218.400 291.000 219.000 ;
        RECT 245.400 217.800 291.000 218.400 ;
        RECT 244.800 217.200 291.000 217.800 ;
        RECT 243.600 216.600 291.000 217.200 ;
        RECT 243.000 216.000 290.400 216.600 ;
        RECT 242.400 215.400 290.400 216.000 ;
        RECT 241.200 214.800 290.400 215.400 ;
        RECT 240.600 214.200 290.400 214.800 ;
        RECT 240.000 213.600 289.800 214.200 ;
        RECT 239.400 213.000 289.800 213.600 ;
        RECT 238.800 212.400 289.800 213.000 ;
        RECT 237.600 211.800 289.800 212.400 ;
        RECT 237.000 211.200 289.200 211.800 ;
        RECT 236.400 210.600 289.200 211.200 ;
        RECT 235.800 210.000 288.600 210.600 ;
        RECT 234.600 209.400 288.600 210.000 ;
        RECT 234.000 208.800 288.000 209.400 ;
        RECT 233.400 208.200 288.000 208.800 ;
        RECT 232.800 207.600 288.000 208.200 ;
        RECT 231.600 207.000 287.400 207.600 ;
        RECT 231.000 206.400 287.400 207.000 ;
        RECT 230.400 205.800 286.800 206.400 ;
        RECT 229.800 205.200 286.800 205.800 ;
        RECT 229.200 204.600 286.200 205.200 ;
        RECT 228.000 204.000 286.200 204.600 ;
        RECT 227.400 203.400 286.200 204.000 ;
        RECT 226.800 202.800 285.600 203.400 ;
        RECT 226.200 202.200 285.600 202.800 ;
        RECT 225.600 201.600 285.000 202.200 ;
        RECT 225.000 201.000 284.400 201.600 ;
        RECT 223.800 200.400 284.400 201.000 ;
        RECT 223.200 199.800 283.800 200.400 ;
        RECT 222.600 199.200 283.800 199.800 ;
        RECT 222.000 198.600 283.200 199.200 ;
        RECT 221.400 198.000 282.600 198.600 ;
        RECT 220.200 197.400 282.600 198.000 ;
        RECT 219.600 196.800 282.000 197.400 ;
        RECT 219.000 196.200 282.000 196.800 ;
        RECT 218.400 195.600 281.400 196.200 ;
        RECT 217.800 195.000 280.800 195.600 ;
        RECT 217.200 194.400 280.800 195.000 ;
        RECT 216.600 193.800 280.200 194.400 ;
        RECT 216.000 193.200 280.200 193.800 ;
        RECT 214.800 192.600 279.600 193.200 ;
        RECT 214.200 192.000 279.000 192.600 ;
        RECT 213.600 191.400 279.000 192.000 ;
        RECT 213.000 190.800 278.400 191.400 ;
        RECT 212.400 190.200 277.800 190.800 ;
        RECT 211.800 189.600 277.800 190.200 ;
        RECT 211.200 189.000 277.200 189.600 ;
        RECT 210.600 188.400 276.600 189.000 ;
        RECT 209.400 187.800 276.000 188.400 ;
        RECT 208.800 187.200 276.000 187.800 ;
        RECT 208.200 186.600 275.400 187.200 ;
        RECT 207.600 186.000 274.800 186.600 ;
        RECT 207.000 185.400 274.800 186.000 ;
        RECT 206.400 184.800 274.200 185.400 ;
        RECT 205.800 184.200 273.600 184.800 ;
        RECT 205.200 183.600 273.000 184.200 ;
        RECT 204.600 183.000 273.000 183.600 ;
        RECT 204.000 182.400 272.400 183.000 ;
        RECT 203.400 181.800 271.800 182.400 ;
        RECT 202.200 181.200 271.800 181.800 ;
        RECT 201.600 180.600 271.200 181.200 ;
        RECT 201.000 180.000 270.600 180.600 ;
        RECT 200.400 179.400 270.000 180.000 ;
        RECT 199.800 178.800 269.400 179.400 ;
        RECT 199.200 178.200 269.400 178.800 ;
        RECT 198.600 177.600 268.800 178.200 ;
        RECT 198.000 177.000 268.200 177.600 ;
        RECT 197.400 176.400 267.600 177.000 ;
        RECT 196.800 175.800 267.600 176.400 ;
        RECT 196.200 175.200 267.000 175.800 ;
        RECT 195.600 174.600 266.400 175.200 ;
        RECT 195.000 174.000 265.800 174.600 ;
        RECT 194.400 173.400 265.200 174.000 ;
        RECT 193.800 172.800 265.200 173.400 ;
        RECT 193.200 172.200 264.600 172.800 ;
        RECT 192.600 171.600 264.000 172.200 ;
        RECT 192.000 171.000 263.400 171.600 ;
        RECT 190.800 170.400 263.400 171.000 ;
        RECT 190.200 169.800 262.800 170.400 ;
        RECT 189.600 169.200 262.200 169.800 ;
        RECT 189.000 168.600 261.600 169.200 ;
        RECT 188.400 168.000 261.000 168.600 ;
        RECT 187.800 167.400 261.000 168.000 ;
        RECT 187.200 166.800 260.400 167.400 ;
        RECT 186.600 166.200 259.800 166.800 ;
        RECT 186.000 165.600 259.200 166.200 ;
        RECT 185.400 165.000 258.600 165.600 ;
        RECT 184.800 164.400 258.600 165.000 ;
        RECT 184.200 163.800 258.000 164.400 ;
        RECT 183.600 163.200 257.400 163.800 ;
        RECT 183.000 162.600 256.800 163.200 ;
        RECT 182.400 162.000 256.200 162.600 ;
        RECT 181.800 161.400 256.200 162.000 ;
        RECT 181.200 160.800 255.600 161.400 ;
        RECT 180.600 160.200 255.000 160.800 ;
        RECT 180.000 159.600 254.400 160.200 ;
        RECT 179.400 159.000 253.800 159.600 ;
        RECT 178.800 158.400 253.200 159.000 ;
        RECT 178.200 157.800 253.200 158.400 ;
        RECT 177.600 157.200 252.600 157.800 ;
        RECT 177.000 156.600 252.000 157.200 ;
        RECT 176.400 156.000 251.400 156.600 ;
        RECT 175.800 155.400 250.800 156.000 ;
        RECT 175.200 154.800 250.800 155.400 ;
        RECT 174.600 154.200 250.200 154.800 ;
        RECT 174.000 153.600 249.600 154.200 ;
        RECT 173.400 153.000 249.000 153.600 ;
        RECT 173.400 152.400 248.400 153.000 ;
        RECT 172.800 151.800 248.400 152.400 ;
        RECT 172.200 151.200 247.800 151.800 ;
        RECT 171.600 150.600 247.200 151.200 ;
        RECT 171.000 150.000 246.600 150.600 ;
        RECT 170.400 149.400 246.000 150.000 ;
        RECT 169.800 148.800 246.000 149.400 ;
        RECT 169.200 148.200 245.400 148.800 ;
        RECT 168.600 147.600 244.800 148.200 ;
        RECT 168.000 147.000 244.200 147.600 ;
        RECT 167.400 146.400 243.600 147.000 ;
        RECT 166.800 145.800 243.000 146.400 ;
        RECT 166.200 145.200 243.000 145.800 ;
        RECT 165.600 144.600 242.400 145.200 ;
        RECT 165.000 144.000 241.800 144.600 ;
        RECT 165.000 143.400 241.200 144.000 ;
        RECT 164.400 142.800 240.600 143.400 ;
        RECT 163.800 142.200 240.600 142.800 ;
        RECT 163.200 141.600 240.000 142.200 ;
        RECT 162.600 141.000 239.400 141.600 ;
        RECT 162.000 140.400 238.800 141.000 ;
        RECT 161.400 139.800 238.200 140.400 ;
        RECT 160.800 139.200 238.200 139.800 ;
        RECT 160.200 138.600 237.600 139.200 ;
        RECT 160.200 138.000 237.000 138.600 ;
        RECT 159.600 137.400 236.400 138.000 ;
        RECT 159.000 136.800 235.800 137.400 ;
        RECT 158.400 136.200 235.200 136.800 ;
        RECT 157.800 135.600 235.200 136.200 ;
        RECT 241.200 135.600 241.800 136.200 ;
        RECT 157.200 135.000 234.600 135.600 ;
        RECT 240.600 135.000 241.800 135.600 ;
        RECT 157.200 134.400 234.000 135.000 ;
        RECT 240.000 134.400 242.400 135.000 ;
        RECT 156.600 133.800 233.400 134.400 ;
        RECT 239.400 133.800 242.400 134.400 ;
        RECT 156.000 133.200 232.800 133.800 ;
        RECT 238.800 133.200 242.400 133.800 ;
        RECT 155.400 132.600 232.800 133.200 ;
        RECT 154.800 132.000 232.200 132.600 ;
        RECT 238.200 132.000 242.400 133.200 ;
        RECT 154.200 131.400 231.600 132.000 ;
        RECT 237.600 131.400 242.400 132.000 ;
        RECT 154.200 130.800 231.000 131.400 ;
        RECT 237.000 130.800 243.000 131.400 ;
        RECT 153.600 130.200 230.400 130.800 ;
        RECT 236.400 130.200 243.000 130.800 ;
        RECT 153.000 129.600 229.800 130.200 ;
        RECT 235.800 129.600 243.000 130.200 ;
        RECT 152.400 129.000 229.800 129.600 ;
        RECT 235.200 129.000 243.000 129.600 ;
        RECT 151.800 128.400 229.200 129.000 ;
        RECT 151.800 127.800 228.600 128.400 ;
        RECT 234.600 127.800 243.000 129.000 ;
        RECT 151.200 127.200 228.000 127.800 ;
        RECT 234.000 127.200 243.000 127.800 ;
        RECT 150.600 126.600 227.400 127.200 ;
        RECT 233.400 126.600 243.000 127.200 ;
        RECT 150.000 126.000 227.400 126.600 ;
        RECT 232.800 126.000 243.000 126.600 ;
        RECT 150.000 125.400 226.800 126.000 ;
        RECT 232.200 125.400 243.000 126.000 ;
        RECT 149.400 124.800 226.200 125.400 ;
        RECT 231.600 124.800 243.000 125.400 ;
        RECT 148.800 124.200 225.600 124.800 ;
        RECT 231.000 124.200 243.000 124.800 ;
        RECT 148.200 123.600 225.000 124.200 ;
        RECT 147.600 123.000 225.000 123.600 ;
        RECT 230.400 123.000 243.000 124.200 ;
        RECT 147.600 122.400 224.400 123.000 ;
        RECT 229.800 122.400 243.000 123.000 ;
        RECT 147.000 121.800 223.800 122.400 ;
        RECT 229.200 121.800 243.000 122.400 ;
        RECT 146.400 121.200 223.200 121.800 ;
        RECT 228.600 121.200 243.000 121.800 ;
        RECT 145.800 120.600 222.600 121.200 ;
        RECT 228.000 120.600 243.000 121.200 ;
        RECT 145.800 120.000 222.000 120.600 ;
        RECT 227.400 120.000 243.000 120.600 ;
        RECT 145.200 119.400 222.000 120.000 ;
        RECT 226.800 119.400 243.000 120.000 ;
        RECT 297.600 119.400 300.000 120.000 ;
        RECT 144.600 118.800 221.400 119.400 ;
        RECT 144.600 118.200 220.800 118.800 ;
        RECT 226.200 118.200 243.000 119.400 ;
        RECT 295.200 118.800 299.400 119.400 ;
        RECT 292.800 118.200 299.400 118.800 ;
        RECT 144.000 117.600 220.200 118.200 ;
        RECT 225.600 117.600 243.000 118.200 ;
        RECT 290.400 117.600 298.800 118.200 ;
        RECT 143.400 117.000 219.600 117.600 ;
        RECT 225.000 117.000 243.000 117.600 ;
        RECT 287.400 117.000 298.800 117.600 ;
        RECT 142.800 116.400 219.600 117.000 ;
        RECT 224.400 116.400 243.000 117.000 ;
        RECT 285.000 116.400 298.800 117.000 ;
        RECT 142.800 115.800 219.000 116.400 ;
        RECT 223.800 115.800 243.000 116.400 ;
        RECT 282.600 115.800 298.200 116.400 ;
        RECT 142.200 115.200 218.400 115.800 ;
        RECT 223.200 115.200 243.000 115.800 ;
        RECT 280.200 115.200 298.200 115.800 ;
        RECT 141.600 114.600 217.800 115.200 ;
        RECT 222.600 114.600 243.000 115.200 ;
        RECT 277.800 114.600 297.600 115.200 ;
        RECT 141.000 114.000 217.200 114.600 ;
        RECT 222.600 114.000 242.400 114.600 ;
        RECT 275.400 114.000 297.600 114.600 ;
        RECT 141.000 113.400 216.600 114.000 ;
        RECT 222.000 113.400 242.400 114.000 ;
        RECT 273.000 113.400 297.600 114.000 ;
        RECT 140.400 112.800 216.600 113.400 ;
        RECT 221.400 112.800 242.400 113.400 ;
        RECT 270.600 112.800 297.000 113.400 ;
        RECT 139.800 112.200 216.000 112.800 ;
        RECT 220.800 112.200 242.400 112.800 ;
        RECT 268.200 112.200 297.000 112.800 ;
        RECT 139.800 111.600 215.400 112.200 ;
        RECT 220.800 111.600 241.200 112.200 ;
        RECT 265.800 111.600 296.400 112.200 ;
        RECT 139.200 111.000 214.800 111.600 ;
        RECT 220.800 111.000 239.400 111.600 ;
        RECT 263.400 111.000 296.400 111.600 ;
        RECT 138.600 109.800 214.200 111.000 ;
        RECT 220.800 110.400 238.200 111.000 ;
        RECT 261.000 110.400 295.800 111.000 ;
        RECT 220.800 109.800 236.400 110.400 ;
        RECT 259.200 109.800 295.800 110.400 ;
        RECT 138.000 109.200 213.600 109.800 ;
        RECT 220.800 109.200 234.600 109.800 ;
        RECT 256.800 109.200 295.200 109.800 ;
        RECT 137.400 108.600 213.000 109.200 ;
        RECT 220.800 108.600 233.400 109.200 ;
        RECT 254.400 108.600 295.200 109.200 ;
        RECT 136.800 108.000 212.400 108.600 ;
        RECT 220.800 108.000 231.600 108.600 ;
        RECT 252.000 108.000 294.600 108.600 ;
        RECT 136.800 107.400 211.800 108.000 ;
        RECT 220.800 107.400 229.800 108.000 ;
        RECT 250.200 107.400 294.600 108.000 ;
        RECT 136.200 106.800 211.200 107.400 ;
        RECT 135.600 106.200 211.200 106.800 ;
        RECT 220.800 106.800 228.000 107.400 ;
        RECT 247.800 106.800 294.000 107.400 ;
        RECT 220.800 106.200 226.800 106.800 ;
        RECT 245.400 106.200 294.000 106.800 ;
        RECT 135.600 105.600 210.600 106.200 ;
        RECT 220.800 105.600 225.000 106.200 ;
        RECT 243.600 105.600 293.400 106.200 ;
        RECT 135.000 105.000 210.000 105.600 ;
        RECT 220.800 105.000 223.200 105.600 ;
        RECT 241.200 105.000 293.400 105.600 ;
        RECT 134.400 104.400 209.400 105.000 ;
        RECT 220.200 104.400 221.400 105.000 ;
        RECT 239.400 104.400 292.800 105.000 ;
        RECT 134.400 103.800 208.800 104.400 ;
        RECT 237.000 103.800 292.200 104.400 ;
        RECT 133.800 103.200 208.200 103.800 ;
        RECT 235.200 103.200 292.200 103.800 ;
        RECT 133.200 102.600 207.000 103.200 ;
        RECT 232.800 102.600 291.600 103.200 ;
        RECT 133.200 102.000 205.800 102.600 ;
        RECT 231.000 102.000 291.600 102.600 ;
        RECT 132.600 101.400 204.600 102.000 ;
        RECT 228.600 101.400 291.000 102.000 ;
        RECT 132.000 100.800 203.400 101.400 ;
        RECT 226.800 100.800 290.400 101.400 ;
        RECT 132.000 100.200 202.200 100.800 ;
        RECT 225.000 100.200 289.800 100.800 ;
        RECT 131.400 99.600 201.000 100.200 ;
        RECT 223.200 99.600 289.200 100.200 ;
        RECT 130.800 99.000 199.800 99.600 ;
        RECT 221.400 99.000 289.200 99.600 ;
        RECT 130.800 98.400 198.600 99.000 ;
        RECT 219.600 98.400 288.600 99.000 ;
        RECT 130.200 97.800 197.400 98.400 ;
        RECT 217.800 97.800 288.000 98.400 ;
        RECT 129.600 97.200 196.200 97.800 ;
        RECT 216.000 97.200 287.400 97.800 ;
        RECT 129.600 96.600 195.000 97.200 ;
        RECT 214.200 96.600 286.800 97.200 ;
        RECT 129.000 96.000 193.800 96.600 ;
        RECT 212.400 96.000 286.200 96.600 ;
        RECT 128.400 95.400 192.600 96.000 ;
        RECT 210.600 95.400 286.200 96.000 ;
        RECT 128.400 94.800 192.000 95.400 ;
        RECT 209.400 94.800 285.600 95.400 ;
        RECT 127.800 94.200 190.800 94.800 ;
        RECT 207.600 94.200 285.000 94.800 ;
        RECT 127.200 93.600 189.600 94.200 ;
        RECT 205.800 93.600 284.400 94.200 ;
        RECT 127.200 93.000 188.400 93.600 ;
        RECT 204.600 93.000 283.800 93.600 ;
        RECT 126.600 92.400 187.200 93.000 ;
        RECT 202.800 92.400 283.200 93.000 ;
        RECT 126.000 91.800 186.000 92.400 ;
        RECT 201.600 91.800 282.600 92.400 ;
        RECT 126.000 91.200 184.800 91.800 ;
        RECT 199.800 91.200 282.000 91.800 ;
        RECT 125.400 90.600 183.600 91.200 ;
        RECT 198.600 90.600 280.800 91.200 ;
        RECT 124.800 90.000 183.000 90.600 ;
        RECT 196.800 90.000 280.200 90.600 ;
        RECT 124.800 89.400 181.800 90.000 ;
        RECT 195.600 89.400 279.600 90.000 ;
        RECT 124.200 88.800 180.600 89.400 ;
        RECT 194.400 88.800 279.000 89.400 ;
        RECT 123.600 88.200 179.400 88.800 ;
        RECT 193.200 88.200 278.400 88.800 ;
        RECT 123.600 87.600 178.200 88.200 ;
        RECT 192.000 87.600 277.200 88.200 ;
        RECT 123.000 87.000 177.000 87.600 ;
        RECT 190.200 87.000 276.600 87.600 ;
        RECT 122.400 86.400 176.400 87.000 ;
        RECT 189.000 86.400 276.000 87.000 ;
        RECT 122.400 85.800 175.200 86.400 ;
        RECT 187.800 85.800 275.400 86.400 ;
        RECT 121.800 85.200 174.000 85.800 ;
        RECT 186.600 85.200 274.200 85.800 ;
        RECT 121.800 84.600 172.800 85.200 ;
        RECT 185.400 84.600 273.600 85.200 ;
        RECT 121.200 84.000 171.600 84.600 ;
        RECT 184.200 84.000 273.000 84.600 ;
        RECT 120.600 83.400 171.000 84.000 ;
        RECT 183.000 83.400 271.800 84.000 ;
        RECT 120.600 82.800 169.800 83.400 ;
        RECT 181.800 82.800 271.200 83.400 ;
        RECT 120.000 82.200 168.600 82.800 ;
        RECT 180.600 82.200 270.000 82.800 ;
        RECT 119.400 81.600 167.400 82.200 ;
        RECT 180.000 81.600 269.400 82.200 ;
        RECT 119.400 81.000 166.800 81.600 ;
        RECT 178.800 81.000 268.800 81.600 ;
        RECT 118.800 80.400 165.600 81.000 ;
        RECT 177.600 80.400 267.600 81.000 ;
        RECT 118.200 79.800 164.400 80.400 ;
        RECT 176.400 79.800 267.000 80.400 ;
        RECT 118.200 79.200 163.800 79.800 ;
        RECT 175.800 79.200 265.800 79.800 ;
        RECT 117.600 78.600 162.600 79.200 ;
        RECT 174.600 78.600 265.200 79.200 ;
        RECT 117.600 78.000 161.400 78.600 ;
        RECT 173.400 78.000 264.000 78.600 ;
        RECT 117.000 77.400 160.800 78.000 ;
        RECT 172.200 77.400 263.400 78.000 ;
        RECT 116.400 76.800 159.600 77.400 ;
        RECT 171.600 76.800 262.200 77.400 ;
        RECT 116.400 76.200 158.400 76.800 ;
        RECT 170.400 76.200 261.000 76.800 ;
        RECT 115.800 75.600 157.800 76.200 ;
        RECT 169.800 75.600 260.400 76.200 ;
        RECT 115.200 75.000 156.600 75.600 ;
        RECT 168.600 75.000 259.200 75.600 ;
        RECT 115.200 74.400 156.000 75.000 ;
        RECT 167.400 74.400 258.600 75.000 ;
        RECT 114.600 73.800 154.800 74.400 ;
        RECT 166.800 73.800 257.400 74.400 ;
        RECT 114.600 73.200 153.600 73.800 ;
        RECT 165.600 73.200 256.800 73.800 ;
        RECT 114.000 72.600 153.000 73.200 ;
        RECT 165.000 72.600 255.600 73.200 ;
        RECT 113.400 72.000 151.800 72.600 ;
        RECT 163.800 72.000 255.000 72.600 ;
        RECT 113.400 71.400 151.200 72.000 ;
        RECT 162.600 71.400 253.800 72.000 ;
        RECT 112.800 70.800 150.000 71.400 ;
        RECT 162.000 70.800 252.600 71.400 ;
        RECT 112.800 70.200 148.800 70.800 ;
        RECT 160.800 70.200 252.000 70.800 ;
        RECT 112.200 69.600 148.200 70.200 ;
        RECT 160.200 69.600 250.800 70.200 ;
        RECT 111.600 69.000 147.000 69.600 ;
        RECT 159.000 69.000 249.600 69.600 ;
        RECT 111.600 68.400 146.400 69.000 ;
        RECT 158.400 68.400 249.000 69.000 ;
        RECT 111.000 67.800 145.200 68.400 ;
        RECT 157.200 67.800 247.800 68.400 ;
        RECT 110.400 67.200 144.600 67.800 ;
        RECT 156.600 67.200 246.600 67.800 ;
        RECT 110.400 66.600 143.400 67.200 ;
        RECT 155.400 66.600 246.000 67.200 ;
        RECT 109.800 66.000 142.800 66.600 ;
        RECT 154.800 66.000 244.800 66.600 ;
        RECT 109.800 65.400 141.600 66.000 ;
        RECT 153.600 65.400 243.600 66.000 ;
        RECT 109.200 64.800 141.000 65.400 ;
        RECT 153.000 64.800 243.000 65.400 ;
        RECT 108.600 64.200 139.800 64.800 ;
        RECT 151.800 64.200 241.800 64.800 ;
        RECT 108.600 63.600 139.200 64.200 ;
        RECT 151.200 63.600 240.600 64.200 ;
        RECT 108.000 63.000 138.000 63.600 ;
        RECT 150.000 63.000 240.000 63.600 ;
        RECT 108.000 62.400 137.400 63.000 ;
        RECT 149.400 62.400 238.800 63.000 ;
        RECT 107.400 61.800 136.800 62.400 ;
        RECT 148.200 61.800 237.600 62.400 ;
        RECT 107.400 61.200 135.600 61.800 ;
        RECT 147.600 61.200 237.000 61.800 ;
        RECT 106.800 60.600 135.000 61.200 ;
        RECT 146.400 60.600 235.800 61.200 ;
        RECT 106.200 60.000 133.800 60.600 ;
        RECT 145.800 60.000 234.600 60.600 ;
        RECT 106.200 59.400 133.200 60.000 ;
        RECT 144.600 59.400 234.000 60.000 ;
        RECT 105.600 58.800 132.000 59.400 ;
        RECT 144.000 58.800 232.800 59.400 ;
        RECT 105.600 58.200 131.400 58.800 ;
        RECT 142.800 58.200 231.600 58.800 ;
        RECT 105.000 57.600 130.800 58.200 ;
        RECT 142.200 57.600 231.000 58.200 ;
        RECT 104.400 57.000 129.600 57.600 ;
        RECT 141.000 57.000 229.800 57.600 ;
        RECT 104.400 56.400 129.000 57.000 ;
        RECT 140.400 56.400 228.600 57.000 ;
        RECT 103.800 55.800 127.800 56.400 ;
        RECT 139.200 55.800 228.000 56.400 ;
        RECT 103.800 55.200 127.200 55.800 ;
        RECT 138.600 55.200 226.800 55.800 ;
        RECT 103.200 54.600 126.600 55.200 ;
        RECT 137.400 54.600 225.600 55.200 ;
        RECT 103.200 54.000 125.400 54.600 ;
        RECT 136.800 54.000 225.000 54.600 ;
        RECT 102.600 53.400 124.800 54.000 ;
        RECT 135.600 53.400 223.800 54.000 ;
        RECT 102.600 52.800 124.200 53.400 ;
        RECT 135.000 52.800 222.600 53.400 ;
        RECT 102.000 52.200 123.000 52.800 ;
        RECT 133.800 52.200 222.000 52.800 ;
        RECT 102.000 51.600 122.400 52.200 ;
        RECT 133.200 51.600 220.800 52.200 ;
        RECT 101.400 51.000 121.800 51.600 ;
        RECT 132.000 51.000 219.600 51.600 ;
        RECT 100.800 50.400 120.600 51.000 ;
        RECT 131.400 50.400 219.000 51.000 ;
        RECT 100.800 49.800 120.000 50.400 ;
        RECT 130.200 49.800 217.800 50.400 ;
        RECT 100.200 49.200 119.400 49.800 ;
        RECT 129.600 49.200 216.600 49.800 ;
        RECT 100.200 48.600 118.800 49.200 ;
        RECT 128.400 48.600 216.000 49.200 ;
        RECT 99.600 48.000 117.600 48.600 ;
        RECT 127.800 48.000 214.800 48.600 ;
        RECT 99.600 47.400 117.000 48.000 ;
        RECT 126.600 47.400 214.200 48.000 ;
        RECT 99.000 46.800 116.400 47.400 ;
        RECT 126.000 46.800 213.000 47.400 ;
        RECT 99.000 46.200 115.200 46.800 ;
        RECT 125.400 46.200 211.800 46.800 ;
        RECT 98.400 45.600 114.600 46.200 ;
        RECT 124.200 45.600 210.600 46.200 ;
        RECT 98.400 45.000 114.000 45.600 ;
        RECT 123.600 45.000 209.400 45.600 ;
        RECT 97.800 44.400 113.400 45.000 ;
        RECT 122.400 44.400 207.600 45.000 ;
        RECT 97.800 43.800 112.200 44.400 ;
        RECT 121.800 43.800 206.400 44.400 ;
        RECT 97.200 43.200 111.600 43.800 ;
        RECT 120.600 43.200 204.600 43.800 ;
        RECT 97.200 42.600 111.000 43.200 ;
        RECT 120.000 42.600 203.400 43.200 ;
        RECT 97.200 42.000 110.400 42.600 ;
        RECT 119.400 42.000 201.600 42.600 ;
        RECT 96.600 41.400 109.200 42.000 ;
        RECT 118.200 41.400 199.800 42.000 ;
        RECT 96.600 40.800 108.600 41.400 ;
        RECT 117.600 40.800 198.600 41.400 ;
        RECT 96.000 40.200 108.000 40.800 ;
        RECT 116.400 40.200 196.800 40.800 ;
        RECT 210.000 40.200 211.200 40.800 ;
        RECT 96.000 39.600 107.400 40.200 ;
        RECT 115.800 39.600 195.600 40.200 ;
        RECT 208.200 39.600 210.600 40.200 ;
        RECT 95.400 39.000 106.200 39.600 ;
        RECT 114.600 39.000 193.800 39.600 ;
        RECT 207.000 39.000 210.000 39.600 ;
        RECT 95.400 38.400 105.600 39.000 ;
        RECT 114.000 38.400 192.600 39.000 ;
        RECT 205.200 38.400 209.400 39.000 ;
        RECT 95.400 37.800 105.000 38.400 ;
        RECT 113.400 37.800 190.800 38.400 ;
        RECT 203.400 37.800 208.800 38.400 ;
        RECT 94.800 37.200 103.800 37.800 ;
        RECT 112.200 37.200 189.600 37.800 ;
        RECT 202.200 37.200 208.200 37.800 ;
        RECT 94.800 36.600 103.200 37.200 ;
        RECT 111.600 36.600 187.800 37.200 ;
        RECT 200.400 36.600 207.600 37.200 ;
        RECT 94.200 36.000 102.600 36.600 ;
        RECT 111.000 36.000 186.600 36.600 ;
        RECT 198.600 36.000 207.000 36.600 ;
        RECT 94.200 35.400 102.000 36.000 ;
        RECT 109.800 35.400 184.800 36.000 ;
        RECT 197.400 35.400 206.400 36.000 ;
        RECT 94.200 34.800 100.800 35.400 ;
        RECT 109.200 34.800 183.600 35.400 ;
        RECT 195.600 34.800 205.200 35.400 ;
        RECT 93.600 34.200 100.200 34.800 ;
        RECT 108.000 34.200 181.800 34.800 ;
        RECT 193.800 34.200 204.600 34.800 ;
        RECT 93.600 33.600 99.600 34.200 ;
        RECT 107.400 33.600 180.000 34.200 ;
        RECT 192.000 33.600 204.000 34.200 ;
        RECT 93.000 33.000 98.400 33.600 ;
        RECT 106.800 33.000 178.800 33.600 ;
        RECT 190.800 33.000 203.400 33.600 ;
        RECT 93.000 32.400 97.800 33.000 ;
        RECT 105.600 32.400 177.000 33.000 ;
        RECT 189.000 32.400 202.800 33.000 ;
        RECT 93.000 31.800 97.200 32.400 ;
        RECT 105.000 31.800 175.800 32.400 ;
        RECT 187.200 31.800 202.200 32.400 ;
        RECT 92.400 31.200 96.000 31.800 ;
        RECT 104.400 31.200 174.000 31.800 ;
        RECT 186.000 31.200 201.600 31.800 ;
        RECT 92.400 30.600 95.400 31.200 ;
        RECT 103.200 30.600 172.800 31.200 ;
        RECT 184.200 30.600 201.000 31.200 ;
        RECT 92.400 30.000 94.800 30.600 ;
        RECT 102.600 30.000 171.000 30.600 ;
        RECT 182.400 30.000 200.400 30.600 ;
        RECT 91.800 29.400 93.600 30.000 ;
        RECT 102.000 29.400 169.800 30.000 ;
        RECT 181.200 29.400 199.800 30.000 ;
        RECT 91.800 28.800 93.000 29.400 ;
        RECT 100.800 28.800 168.000 29.400 ;
        RECT 179.400 28.800 198.600 29.400 ;
        RECT 91.200 28.200 92.400 28.800 ;
        RECT 100.200 28.200 124.200 28.800 ;
        RECT 177.600 28.200 198.000 28.800 ;
        RECT 99.600 27.600 120.000 28.200 ;
        RECT 176.400 27.600 197.400 28.200 ;
        RECT 98.400 27.000 117.600 27.600 ;
        RECT 174.600 27.000 196.800 27.600 ;
        RECT 97.800 26.400 115.200 27.000 ;
        RECT 172.800 26.400 196.200 27.000 ;
        RECT 97.200 25.800 114.000 26.400 ;
        RECT 171.600 25.800 195.600 26.400 ;
        RECT 96.600 25.200 112.200 25.800 ;
        RECT 169.800 25.200 195.000 25.800 ;
        RECT 96.000 24.600 111.000 25.200 ;
        RECT 150.600 24.600 193.800 25.200 ;
        RECT 94.800 24.000 109.800 24.600 ;
        RECT 148.200 24.000 193.200 24.600 ;
        RECT 94.200 23.400 108.000 24.000 ;
        RECT 146.400 23.400 192.600 24.000 ;
        RECT 93.600 22.800 107.400 23.400 ;
        RECT 144.000 22.800 191.400 23.400 ;
        RECT 93.000 22.200 106.200 22.800 ;
        RECT 141.000 22.200 190.800 22.800 ;
        RECT 92.400 21.600 105.000 22.200 ;
        RECT 137.400 21.600 190.200 22.200 ;
        RECT 91.800 21.000 103.800 21.600 ;
        RECT 132.600 21.000 189.600 21.600 ;
        RECT 91.200 20.400 103.200 21.000 ;
        RECT 109.200 20.400 117.000 21.000 ;
        RECT 124.200 20.400 188.400 21.000 ;
        RECT 90.600 19.800 102.000 20.400 ;
        RECT 108.600 19.800 187.800 20.400 ;
        RECT 90.000 19.200 101.400 19.800 ;
        RECT 108.000 19.200 186.600 19.800 ;
        RECT 89.400 18.600 100.200 19.200 ;
        RECT 106.800 18.600 186.000 19.200 ;
        RECT 88.800 18.000 99.600 18.600 ;
        RECT 106.200 18.000 184.800 18.600 ;
        RECT 88.200 17.400 98.400 18.000 ;
        RECT 105.600 17.400 184.200 18.000 ;
        RECT 88.200 16.800 97.800 17.400 ;
        RECT 105.000 16.800 183.000 17.400 ;
        RECT 87.600 16.200 97.200 16.800 ;
        RECT 104.400 16.200 182.400 16.800 ;
        RECT 87.000 15.600 96.000 16.200 ;
        RECT 103.200 15.600 181.200 16.200 ;
        RECT 87.000 15.000 95.400 15.600 ;
        RECT 102.600 15.000 180.000 15.600 ;
        RECT 86.400 14.400 94.800 15.000 ;
        RECT 102.000 14.400 179.400 15.000 ;
        RECT 85.800 13.800 93.600 14.400 ;
        RECT 101.400 13.800 178.200 14.400 ;
        RECT 85.800 13.200 93.000 13.800 ;
        RECT 100.200 13.200 177.000 13.800 ;
        RECT 85.200 12.600 92.400 13.200 ;
        RECT 99.600 12.600 175.800 13.200 ;
        RECT 85.200 12.000 91.200 12.600 ;
        RECT 99.000 12.000 174.600 12.600 ;
        RECT 84.600 11.400 90.600 12.000 ;
        RECT 98.400 11.400 173.400 12.000 ;
        RECT 84.600 10.800 89.400 11.400 ;
        RECT 97.200 10.800 172.200 11.400 ;
        RECT 84.000 10.200 88.800 10.800 ;
        RECT 96.600 10.200 171.000 10.800 ;
        RECT 84.000 9.600 87.600 10.200 ;
        RECT 96.000 9.600 169.800 10.200 ;
        RECT 83.400 9.000 87.000 9.600 ;
        RECT 95.400 9.000 168.000 9.600 ;
        RECT 83.400 8.400 85.800 9.000 ;
        RECT 94.800 8.400 166.800 9.000 ;
        RECT 82.800 7.800 84.600 8.400 ;
        RECT 93.600 7.800 165.000 8.400 ;
        RECT 82.800 7.200 84.000 7.800 ;
        RECT 93.000 7.200 163.800 7.800 ;
        RECT 92.400 6.600 162.000 7.200 ;
        RECT 91.800 6.000 160.200 6.600 ;
        RECT 90.600 5.400 158.400 6.000 ;
        RECT 90.000 4.800 156.600 5.400 ;
        RECT 89.400 4.200 154.200 4.800 ;
        RECT 91.800 3.600 152.400 4.200 ;
        RECT 95.400 3.000 150.000 3.600 ;
        RECT 99.600 2.400 147.000 3.000 ;
        RECT 103.200 1.800 144.600 2.400 ;
        RECT 108.000 1.200 141.000 1.800 ;
        RECT 112.800 0.600 136.800 1.200 ;
        RECT 121.200 0.000 128.400 0.600 ;
  END
END avali_logo
END LIBRARY

