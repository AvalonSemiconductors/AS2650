// This is the unpowered netlist.
module wrapped_as2650 (WEb_raw,
    boot_rom_en,
    bus_cyc,
    bus_we_gpios,
    bus_we_serial_ports,
    bus_we_timers,
    le_hi_act,
    le_lo_act,
    reset_out,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    RAM_end_addr,
    RAM_start_addr,
    bus_addr,
    bus_data_out,
    bus_in_gpios,
    bus_in_serial_ports,
    bus_in_timers,
    cs_port,
    io_in,
    io_oeb,
    io_out,
    irq,
    irqs,
    la_data_out,
    rom_bus_in,
    rom_bus_out,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o);
 output WEb_raw;
 output boot_rom_en;
 output bus_cyc;
 output bus_we_gpios;
 output bus_we_serial_ports;
 output bus_we_timers;
 output le_hi_act;
 output le_lo_act;
 output reset_out;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 output [15:0] RAM_end_addr;
 output [15:0] RAM_start_addr;
 output [5:0] bus_addr;
 output [7:0] bus_data_out;
 input [7:0] bus_in_gpios;
 input [7:0] bus_in_serial_ports;
 input [7:0] bus_in_timers;
 output [2:0] cs_port;
 input [18:0] io_in;
 output [18:0] io_oeb;
 output [18:0] io_out;
 output [2:0] irq;
 input [6:0] irqs;
 output [55:0] la_data_out;
 input [7:0] rom_bus_in;
 output [7:0] rom_bus_out;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;

 wire net275;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net254;
 wire net255;
 wire net276;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire \as2650.PC[0] ;
 wire \as2650.PC[10] ;
 wire \as2650.PC[11] ;
 wire \as2650.PC[12] ;
 wire \as2650.PC[1] ;
 wire \as2650.PC[2] ;
 wire \as2650.PC[3] ;
 wire \as2650.PC[4] ;
 wire \as2650.PC[5] ;
 wire \as2650.PC[6] ;
 wire \as2650.PC[7] ;
 wire \as2650.PC[8] ;
 wire \as2650.PC[9] ;
 wire \as2650.chirp_ptr[0] ;
 wire \as2650.chirp_ptr[1] ;
 wire \as2650.chirp_ptr[2] ;
 wire \as2650.chirpchar[0] ;
 wire \as2650.chirpchar[1] ;
 wire \as2650.chirpchar[2] ;
 wire \as2650.chirpchar[3] ;
 wire \as2650.chirpchar[4] ;
 wire \as2650.chirpchar[5] ;
 wire \as2650.chirpchar[6] ;
 wire \as2650.cpu_hidden_rom_enable ;
 wire \as2650.cycle[0] ;
 wire \as2650.cycle[1] ;
 wire \as2650.cycle[2] ;
 wire \as2650.cycle[3] ;
 wire \as2650.debug_psl[0] ;
 wire \as2650.debug_psl[1] ;
 wire \as2650.debug_psl[2] ;
 wire \as2650.debug_psl[3] ;
 wire \as2650.debug_psl[4] ;
 wire \as2650.debug_psl[5] ;
 wire \as2650.debug_psl[6] ;
 wire \as2650.debug_psl[7] ;
 wire \as2650.debug_psu[0] ;
 wire \as2650.debug_psu[1] ;
 wire \as2650.debug_psu[2] ;
 wire \as2650.debug_psu[3] ;
 wire \as2650.debug_psu[4] ;
 wire \as2650.debug_psu[5] ;
 wire \as2650.debug_psu[7] ;
 wire \as2650.ext_io_addr[6] ;
 wire \as2650.ext_io_addr[7] ;
 wire \as2650.extend ;
 wire \as2650.indexed_cyc[0] ;
 wire \as2650.indexed_cyc[1] ;
 wire \as2650.indirect_cyc ;
 wire \as2650.indirect_target[0] ;
 wire \as2650.indirect_target[10] ;
 wire \as2650.indirect_target[11] ;
 wire \as2650.indirect_target[12] ;
 wire \as2650.indirect_target[13] ;
 wire \as2650.indirect_target[14] ;
 wire \as2650.indirect_target[15] ;
 wire \as2650.indirect_target[1] ;
 wire \as2650.indirect_target[2] ;
 wire \as2650.indirect_target[3] ;
 wire \as2650.indirect_target[4] ;
 wire \as2650.indirect_target[5] ;
 wire \as2650.indirect_target[6] ;
 wire \as2650.indirect_target[7] ;
 wire \as2650.indirect_target[8] ;
 wire \as2650.indirect_target[9] ;
 wire \as2650.insin[0] ;
 wire \as2650.insin[1] ;
 wire \as2650.insin[2] ;
 wire \as2650.insin[3] ;
 wire \as2650.insin[4] ;
 wire \as2650.insin[5] ;
 wire \as2650.insin[6] ;
 wire \as2650.insin[7] ;
 wire \as2650.instruction_args_latch[0] ;
 wire \as2650.instruction_args_latch[10] ;
 wire \as2650.instruction_args_latch[11] ;
 wire \as2650.instruction_args_latch[12] ;
 wire \as2650.instruction_args_latch[13] ;
 wire \as2650.instruction_args_latch[14] ;
 wire \as2650.instruction_args_latch[15] ;
 wire \as2650.instruction_args_latch[1] ;
 wire \as2650.instruction_args_latch[2] ;
 wire \as2650.instruction_args_latch[3] ;
 wire \as2650.instruction_args_latch[4] ;
 wire \as2650.instruction_args_latch[5] ;
 wire \as2650.instruction_args_latch[6] ;
 wire \as2650.instruction_args_latch[7] ;
 wire \as2650.instruction_args_latch[8] ;
 wire \as2650.instruction_args_latch[9] ;
 wire \as2650.io_bus_we ;
 wire \as2650.irqs_latch[1] ;
 wire \as2650.irqs_latch[2] ;
 wire \as2650.irqs_latch[3] ;
 wire \as2650.irqs_latch[4] ;
 wire \as2650.irqs_latch[5] ;
 wire \as2650.irqs_latch[6] ;
 wire \as2650.irqs_latch[7] ;
 wire \as2650.ivectors_base[0] ;
 wire \as2650.ivectors_base[10] ;
 wire \as2650.ivectors_base[11] ;
 wire \as2650.ivectors_base[1] ;
 wire \as2650.ivectors_base[2] ;
 wire \as2650.ivectors_base[3] ;
 wire \as2650.ivectors_base[4] ;
 wire \as2650.ivectors_base[5] ;
 wire \as2650.ivectors_base[6] ;
 wire \as2650.ivectors_base[7] ;
 wire \as2650.ivectors_base[8] ;
 wire \as2650.ivectors_base[9] ;
 wire \as2650.last_addr[0] ;
 wire \as2650.last_addr[10] ;
 wire \as2650.last_addr[11] ;
 wire \as2650.last_addr[12] ;
 wire \as2650.last_addr[13] ;
 wire \as2650.last_addr[14] ;
 wire \as2650.last_addr[15] ;
 wire \as2650.last_addr[1] ;
 wire \as2650.last_addr[2] ;
 wire \as2650.last_addr[3] ;
 wire \as2650.last_addr[4] ;
 wire \as2650.last_addr[5] ;
 wire \as2650.last_addr[6] ;
 wire \as2650.last_addr[7] ;
 wire \as2650.last_addr[8] ;
 wire \as2650.last_addr[9] ;
 wire \as2650.page_reg[0] ;
 wire \as2650.page_reg[1] ;
 wire \as2650.page_reg[2] ;
 wire \as2650.regs[0][0] ;
 wire \as2650.regs[0][1] ;
 wire \as2650.regs[0][2] ;
 wire \as2650.regs[0][3] ;
 wire \as2650.regs[0][4] ;
 wire \as2650.regs[0][5] ;
 wire \as2650.regs[0][6] ;
 wire \as2650.regs[0][7] ;
 wire \as2650.regs[1][0] ;
 wire \as2650.regs[1][1] ;
 wire \as2650.regs[1][2] ;
 wire \as2650.regs[1][3] ;
 wire \as2650.regs[1][4] ;
 wire \as2650.regs[1][5] ;
 wire \as2650.regs[1][6] ;
 wire \as2650.regs[1][7] ;
 wire \as2650.regs[2][0] ;
 wire \as2650.regs[2][1] ;
 wire \as2650.regs[2][2] ;
 wire \as2650.regs[2][3] ;
 wire \as2650.regs[2][4] ;
 wire \as2650.regs[2][5] ;
 wire \as2650.regs[2][6] ;
 wire \as2650.regs[2][7] ;
 wire \as2650.regs[3][0] ;
 wire \as2650.regs[3][1] ;
 wire \as2650.regs[3][2] ;
 wire \as2650.regs[3][3] ;
 wire \as2650.regs[3][4] ;
 wire \as2650.regs[3][5] ;
 wire \as2650.regs[3][6] ;
 wire \as2650.regs[3][7] ;
 wire \as2650.regs[4][0] ;
 wire \as2650.regs[4][1] ;
 wire \as2650.regs[4][2] ;
 wire \as2650.regs[4][3] ;
 wire \as2650.regs[4][4] ;
 wire \as2650.regs[4][5] ;
 wire \as2650.regs[4][6] ;
 wire \as2650.regs[4][7] ;
 wire \as2650.regs[5][0] ;
 wire \as2650.regs[5][1] ;
 wire \as2650.regs[5][2] ;
 wire \as2650.regs[5][3] ;
 wire \as2650.regs[5][4] ;
 wire \as2650.regs[5][5] ;
 wire \as2650.regs[5][6] ;
 wire \as2650.regs[5][7] ;
 wire \as2650.regs[6][0] ;
 wire \as2650.regs[6][1] ;
 wire \as2650.regs[6][2] ;
 wire \as2650.regs[6][3] ;
 wire \as2650.regs[6][4] ;
 wire \as2650.regs[6][5] ;
 wire \as2650.regs[6][6] ;
 wire \as2650.regs[6][7] ;
 wire \as2650.regs[7][0] ;
 wire \as2650.regs[7][1] ;
 wire \as2650.regs[7][2] ;
 wire \as2650.regs[7][3] ;
 wire \as2650.regs[7][4] ;
 wire \as2650.regs[7][5] ;
 wire \as2650.regs[7][6] ;
 wire \as2650.regs[7][7] ;
 wire \as2650.relative_cyc ;
 wire \as2650.stack[0][0] ;
 wire \as2650.stack[0][10] ;
 wire \as2650.stack[0][11] ;
 wire \as2650.stack[0][12] ;
 wire \as2650.stack[0][13] ;
 wire \as2650.stack[0][14] ;
 wire \as2650.stack[0][15] ;
 wire \as2650.stack[0][1] ;
 wire \as2650.stack[0][2] ;
 wire \as2650.stack[0][3] ;
 wire \as2650.stack[0][4] ;
 wire \as2650.stack[0][5] ;
 wire \as2650.stack[0][6] ;
 wire \as2650.stack[0][7] ;
 wire \as2650.stack[0][8] ;
 wire \as2650.stack[0][9] ;
 wire \as2650.stack[10][0] ;
 wire \as2650.stack[10][10] ;
 wire \as2650.stack[10][11] ;
 wire \as2650.stack[10][12] ;
 wire \as2650.stack[10][13] ;
 wire \as2650.stack[10][14] ;
 wire \as2650.stack[10][15] ;
 wire \as2650.stack[10][1] ;
 wire \as2650.stack[10][2] ;
 wire \as2650.stack[10][3] ;
 wire \as2650.stack[10][4] ;
 wire \as2650.stack[10][5] ;
 wire \as2650.stack[10][6] ;
 wire \as2650.stack[10][7] ;
 wire \as2650.stack[10][8] ;
 wire \as2650.stack[10][9] ;
 wire \as2650.stack[11][0] ;
 wire \as2650.stack[11][10] ;
 wire \as2650.stack[11][11] ;
 wire \as2650.stack[11][12] ;
 wire \as2650.stack[11][13] ;
 wire \as2650.stack[11][14] ;
 wire \as2650.stack[11][15] ;
 wire \as2650.stack[11][1] ;
 wire \as2650.stack[11][2] ;
 wire \as2650.stack[11][3] ;
 wire \as2650.stack[11][4] ;
 wire \as2650.stack[11][5] ;
 wire \as2650.stack[11][6] ;
 wire \as2650.stack[11][7] ;
 wire \as2650.stack[11][8] ;
 wire \as2650.stack[11][9] ;
 wire \as2650.stack[12][0] ;
 wire \as2650.stack[12][10] ;
 wire \as2650.stack[12][11] ;
 wire \as2650.stack[12][12] ;
 wire \as2650.stack[12][13] ;
 wire \as2650.stack[12][14] ;
 wire \as2650.stack[12][15] ;
 wire \as2650.stack[12][1] ;
 wire \as2650.stack[12][2] ;
 wire \as2650.stack[12][3] ;
 wire \as2650.stack[12][4] ;
 wire \as2650.stack[12][5] ;
 wire \as2650.stack[12][6] ;
 wire \as2650.stack[12][7] ;
 wire \as2650.stack[12][8] ;
 wire \as2650.stack[12][9] ;
 wire \as2650.stack[13][0] ;
 wire \as2650.stack[13][10] ;
 wire \as2650.stack[13][11] ;
 wire \as2650.stack[13][12] ;
 wire \as2650.stack[13][13] ;
 wire \as2650.stack[13][14] ;
 wire \as2650.stack[13][15] ;
 wire \as2650.stack[13][1] ;
 wire \as2650.stack[13][2] ;
 wire \as2650.stack[13][3] ;
 wire \as2650.stack[13][4] ;
 wire \as2650.stack[13][5] ;
 wire \as2650.stack[13][6] ;
 wire \as2650.stack[13][7] ;
 wire \as2650.stack[13][8] ;
 wire \as2650.stack[13][9] ;
 wire \as2650.stack[14][0] ;
 wire \as2650.stack[14][10] ;
 wire \as2650.stack[14][11] ;
 wire \as2650.stack[14][12] ;
 wire \as2650.stack[14][13] ;
 wire \as2650.stack[14][14] ;
 wire \as2650.stack[14][15] ;
 wire \as2650.stack[14][1] ;
 wire \as2650.stack[14][2] ;
 wire \as2650.stack[14][3] ;
 wire \as2650.stack[14][4] ;
 wire \as2650.stack[14][5] ;
 wire \as2650.stack[14][6] ;
 wire \as2650.stack[14][7] ;
 wire \as2650.stack[14][8] ;
 wire \as2650.stack[14][9] ;
 wire \as2650.stack[15][0] ;
 wire \as2650.stack[15][10] ;
 wire \as2650.stack[15][11] ;
 wire \as2650.stack[15][12] ;
 wire \as2650.stack[15][13] ;
 wire \as2650.stack[15][14] ;
 wire \as2650.stack[15][15] ;
 wire \as2650.stack[15][1] ;
 wire \as2650.stack[15][2] ;
 wire \as2650.stack[15][3] ;
 wire \as2650.stack[15][4] ;
 wire \as2650.stack[15][5] ;
 wire \as2650.stack[15][6] ;
 wire \as2650.stack[15][7] ;
 wire \as2650.stack[15][8] ;
 wire \as2650.stack[15][9] ;
 wire \as2650.stack[1][0] ;
 wire \as2650.stack[1][10] ;
 wire \as2650.stack[1][11] ;
 wire \as2650.stack[1][12] ;
 wire \as2650.stack[1][13] ;
 wire \as2650.stack[1][14] ;
 wire \as2650.stack[1][15] ;
 wire \as2650.stack[1][1] ;
 wire \as2650.stack[1][2] ;
 wire \as2650.stack[1][3] ;
 wire \as2650.stack[1][4] ;
 wire \as2650.stack[1][5] ;
 wire \as2650.stack[1][6] ;
 wire \as2650.stack[1][7] ;
 wire \as2650.stack[1][8] ;
 wire \as2650.stack[1][9] ;
 wire \as2650.stack[2][0] ;
 wire \as2650.stack[2][10] ;
 wire \as2650.stack[2][11] ;
 wire \as2650.stack[2][12] ;
 wire \as2650.stack[2][13] ;
 wire \as2650.stack[2][14] ;
 wire \as2650.stack[2][15] ;
 wire \as2650.stack[2][1] ;
 wire \as2650.stack[2][2] ;
 wire \as2650.stack[2][3] ;
 wire \as2650.stack[2][4] ;
 wire \as2650.stack[2][5] ;
 wire \as2650.stack[2][6] ;
 wire \as2650.stack[2][7] ;
 wire \as2650.stack[2][8] ;
 wire \as2650.stack[2][9] ;
 wire \as2650.stack[3][0] ;
 wire \as2650.stack[3][10] ;
 wire \as2650.stack[3][11] ;
 wire \as2650.stack[3][12] ;
 wire \as2650.stack[3][13] ;
 wire \as2650.stack[3][14] ;
 wire \as2650.stack[3][15] ;
 wire \as2650.stack[3][1] ;
 wire \as2650.stack[3][2] ;
 wire \as2650.stack[3][3] ;
 wire \as2650.stack[3][4] ;
 wire \as2650.stack[3][5] ;
 wire \as2650.stack[3][6] ;
 wire \as2650.stack[3][7] ;
 wire \as2650.stack[3][8] ;
 wire \as2650.stack[3][9] ;
 wire \as2650.stack[4][0] ;
 wire \as2650.stack[4][10] ;
 wire \as2650.stack[4][11] ;
 wire \as2650.stack[4][12] ;
 wire \as2650.stack[4][13] ;
 wire \as2650.stack[4][14] ;
 wire \as2650.stack[4][15] ;
 wire \as2650.stack[4][1] ;
 wire \as2650.stack[4][2] ;
 wire \as2650.stack[4][3] ;
 wire \as2650.stack[4][4] ;
 wire \as2650.stack[4][5] ;
 wire \as2650.stack[4][6] ;
 wire \as2650.stack[4][7] ;
 wire \as2650.stack[4][8] ;
 wire \as2650.stack[4][9] ;
 wire \as2650.stack[5][0] ;
 wire \as2650.stack[5][10] ;
 wire \as2650.stack[5][11] ;
 wire \as2650.stack[5][12] ;
 wire \as2650.stack[5][13] ;
 wire \as2650.stack[5][14] ;
 wire \as2650.stack[5][15] ;
 wire \as2650.stack[5][1] ;
 wire \as2650.stack[5][2] ;
 wire \as2650.stack[5][3] ;
 wire \as2650.stack[5][4] ;
 wire \as2650.stack[5][5] ;
 wire \as2650.stack[5][6] ;
 wire \as2650.stack[5][7] ;
 wire \as2650.stack[5][8] ;
 wire \as2650.stack[5][9] ;
 wire \as2650.stack[6][0] ;
 wire \as2650.stack[6][10] ;
 wire \as2650.stack[6][11] ;
 wire \as2650.stack[6][12] ;
 wire \as2650.stack[6][13] ;
 wire \as2650.stack[6][14] ;
 wire \as2650.stack[6][15] ;
 wire \as2650.stack[6][1] ;
 wire \as2650.stack[6][2] ;
 wire \as2650.stack[6][3] ;
 wire \as2650.stack[6][4] ;
 wire \as2650.stack[6][5] ;
 wire \as2650.stack[6][6] ;
 wire \as2650.stack[6][7] ;
 wire \as2650.stack[6][8] ;
 wire \as2650.stack[6][9] ;
 wire \as2650.stack[7][0] ;
 wire \as2650.stack[7][10] ;
 wire \as2650.stack[7][11] ;
 wire \as2650.stack[7][12] ;
 wire \as2650.stack[7][13] ;
 wire \as2650.stack[7][14] ;
 wire \as2650.stack[7][15] ;
 wire \as2650.stack[7][1] ;
 wire \as2650.stack[7][2] ;
 wire \as2650.stack[7][3] ;
 wire \as2650.stack[7][4] ;
 wire \as2650.stack[7][5] ;
 wire \as2650.stack[7][6] ;
 wire \as2650.stack[7][7] ;
 wire \as2650.stack[7][8] ;
 wire \as2650.stack[7][9] ;
 wire \as2650.stack[8][0] ;
 wire \as2650.stack[8][10] ;
 wire \as2650.stack[8][11] ;
 wire \as2650.stack[8][12] ;
 wire \as2650.stack[8][13] ;
 wire \as2650.stack[8][14] ;
 wire \as2650.stack[8][15] ;
 wire \as2650.stack[8][1] ;
 wire \as2650.stack[8][2] ;
 wire \as2650.stack[8][3] ;
 wire \as2650.stack[8][4] ;
 wire \as2650.stack[8][5] ;
 wire \as2650.stack[8][6] ;
 wire \as2650.stack[8][7] ;
 wire \as2650.stack[8][8] ;
 wire \as2650.stack[8][9] ;
 wire \as2650.stack[9][0] ;
 wire \as2650.stack[9][10] ;
 wire \as2650.stack[9][11] ;
 wire \as2650.stack[9][12] ;
 wire \as2650.stack[9][13] ;
 wire \as2650.stack[9][14] ;
 wire \as2650.stack[9][15] ;
 wire \as2650.stack[9][1] ;
 wire \as2650.stack[9][2] ;
 wire \as2650.stack[9][3] ;
 wire \as2650.stack[9][4] ;
 wire \as2650.stack[9][5] ;
 wire \as2650.stack[9][6] ;
 wire \as2650.stack[9][7] ;
 wire \as2650.stack[9][8] ;
 wire \as2650.stack[9][9] ;
 wire \as2650.trap ;
 wire \as2650.warmup[0] ;
 wire \as2650.warmup[1] ;
 wire \as2650.wb_hidden_rom_enable ;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_wb_clk_i;
 wire clknet_4_0__leaf_wb_clk_i;
 wire clknet_4_10__leaf_wb_clk_i;
 wire clknet_4_11__leaf_wb_clk_i;
 wire clknet_4_12__leaf_wb_clk_i;
 wire clknet_4_13__leaf_wb_clk_i;
 wire clknet_4_14__leaf_wb_clk_i;
 wire clknet_4_15__leaf_wb_clk_i;
 wire clknet_4_1__leaf_wb_clk_i;
 wire clknet_4_2__leaf_wb_clk_i;
 wire clknet_4_3__leaf_wb_clk_i;
 wire clknet_4_4__leaf_wb_clk_i;
 wire clknet_4_5__leaf_wb_clk_i;
 wire clknet_4_6__leaf_wb_clk_i;
 wire clknet_4_7__leaf_wb_clk_i;
 wire clknet_4_8__leaf_wb_clk_i;
 wire clknet_4_9__leaf_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_101_wb_clk_i;
 wire clknet_leaf_102_wb_clk_i;
 wire clknet_leaf_103_wb_clk_i;
 wire clknet_leaf_104_wb_clk_i;
 wire clknet_leaf_105_wb_clk_i;
 wire clknet_leaf_106_wb_clk_i;
 wire clknet_leaf_107_wb_clk_i;
 wire clknet_leaf_108_wb_clk_i;
 wire clknet_leaf_109_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_110_wb_clk_i;
 wire clknet_leaf_111_wb_clk_i;
 wire clknet_leaf_112_wb_clk_i;
 wire clknet_leaf_113_wb_clk_i;
 wire clknet_leaf_114_wb_clk_i;
 wire clknet_leaf_115_wb_clk_i;
 wire clknet_leaf_116_wb_clk_i;
 wire clknet_leaf_117_wb_clk_i;
 wire clknet_leaf_118_wb_clk_i;
 wire clknet_leaf_119_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_120_wb_clk_i;
 wire clknet_leaf_121_wb_clk_i;
 wire clknet_leaf_122_wb_clk_i;
 wire clknet_leaf_123_wb_clk_i;
 wire clknet_leaf_124_wb_clk_i;
 wire clknet_leaf_125_wb_clk_i;
 wire clknet_leaf_126_wb_clk_i;
 wire clknet_leaf_127_wb_clk_i;
 wire clknet_leaf_128_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_130_wb_clk_i;
 wire clknet_leaf_131_wb_clk_i;
 wire clknet_leaf_132_wb_clk_i;
 wire clknet_leaf_133_wb_clk_i;
 wire clknet_leaf_134_wb_clk_i;
 wire clknet_leaf_135_wb_clk_i;
 wire clknet_leaf_136_wb_clk_i;
 wire clknet_leaf_137_wb_clk_i;
 wire clknet_leaf_138_wb_clk_i;
 wire clknet_leaf_139_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_140_wb_clk_i;
 wire clknet_leaf_141_wb_clk_i;
 wire clknet_leaf_142_wb_clk_i;
 wire clknet_leaf_143_wb_clk_i;
 wire clknet_leaf_144_wb_clk_i;
 wire clknet_leaf_145_wb_clk_i;
 wire clknet_leaf_146_wb_clk_i;
 wire clknet_leaf_147_wb_clk_i;
 wire clknet_leaf_148_wb_clk_i;
 wire clknet_leaf_149_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_150_wb_clk_i;
 wire clknet_leaf_152_wb_clk_i;
 wire clknet_leaf_153_wb_clk_i;
 wire clknet_leaf_154_wb_clk_i;
 wire clknet_leaf_155_wb_clk_i;
 wire clknet_leaf_156_wb_clk_i;
 wire clknet_leaf_157_wb_clk_i;
 wire clknet_leaf_158_wb_clk_i;
 wire clknet_leaf_159_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_160_wb_clk_i;
 wire clknet_leaf_161_wb_clk_i;
 wire clknet_leaf_162_wb_clk_i;
 wire clknet_leaf_163_wb_clk_i;
 wire clknet_leaf_164_wb_clk_i;
 wire clknet_leaf_165_wb_clk_i;
 wire clknet_leaf_166_wb_clk_i;
 wire clknet_leaf_167_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_57_wb_clk_i;
 wire clknet_leaf_58_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_60_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_62_wb_clk_i;
 wire clknet_leaf_64_wb_clk_i;
 wire clknet_leaf_66_wb_clk_i;
 wire clknet_leaf_67_wb_clk_i;
 wire clknet_leaf_68_wb_clk_i;
 wire clknet_leaf_69_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_70_wb_clk_i;
 wire clknet_leaf_71_wb_clk_i;
 wire clknet_leaf_72_wb_clk_i;
 wire clknet_leaf_73_wb_clk_i;
 wire clknet_leaf_74_wb_clk_i;
 wire clknet_leaf_75_wb_clk_i;
 wire clknet_leaf_76_wb_clk_i;
 wire clknet_leaf_77_wb_clk_i;
 wire clknet_leaf_78_wb_clk_i;
 wire clknet_leaf_79_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_80_wb_clk_i;
 wire clknet_leaf_81_wb_clk_i;
 wire clknet_leaf_82_wb_clk_i;
 wire clknet_leaf_83_wb_clk_i;
 wire clknet_leaf_85_wb_clk_i;
 wire clknet_leaf_87_wb_clk_i;
 wire clknet_leaf_88_wb_clk_i;
 wire clknet_leaf_89_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_90_wb_clk_i;
 wire clknet_leaf_91_wb_clk_i;
 wire clknet_leaf_92_wb_clk_i;
 wire clknet_leaf_93_wb_clk_i;
 wire clknet_leaf_94_wb_clk_i;
 wire clknet_leaf_95_wb_clk_i;
 wire clknet_leaf_96_wb_clk_i;
 wire clknet_leaf_97_wb_clk_i;
 wire clknet_leaf_98_wb_clk_i;
 wire clknet_leaf_99_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \wb_counter[0] ;
 wire \wb_counter[10] ;
 wire \wb_counter[11] ;
 wire \wb_counter[12] ;
 wire \wb_counter[13] ;
 wire \wb_counter[14] ;
 wire \wb_counter[15] ;
 wire \wb_counter[16] ;
 wire \wb_counter[17] ;
 wire \wb_counter[18] ;
 wire \wb_counter[19] ;
 wire \wb_counter[1] ;
 wire \wb_counter[20] ;
 wire \wb_counter[21] ;
 wire \wb_counter[22] ;
 wire \wb_counter[23] ;
 wire \wb_counter[24] ;
 wire \wb_counter[25] ;
 wire \wb_counter[26] ;
 wire \wb_counter[27] ;
 wire \wb_counter[28] ;
 wire \wb_counter[29] ;
 wire \wb_counter[2] ;
 wire \wb_counter[30] ;
 wire \wb_counter[31] ;
 wire \wb_counter[3] ;
 wire \wb_counter[4] ;
 wire \wb_counter[5] ;
 wire \wb_counter[6] ;
 wire \wb_counter[7] ;
 wire \wb_counter[8] ;
 wire \wb_counter[9] ;
 wire wb_debug_carry;
 wire wb_debug_cc;
 wire wb_feedback_delay;
 wire wb_io3_test;
 wire wb_reset_override;
 wire wb_reset_override_en;
 wire \web_behavior[0] ;
 wire \web_behavior[1] ;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05743__I0 (.I(\as2650.regs[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05743__I1 (.I(\as2650.regs[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05744__I (.I(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05748__I0 (.I(\as2650.regs[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05748__I1 (.I(\as2650.regs[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05749__I (.I(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05752__S (.I(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05753__I (.I(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05756__I1 (.I(\as2650.regs[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05756__S (.I(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05758__I (.I(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05759__I1 (.I(\as2650.regs[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05760__I (.I(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05763__I0 (.I(\as2650.regs[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05763__I1 (.I(\as2650.regs[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05767__I0 (.I(\as2650.regs[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05767__I1 (.I(\as2650.regs[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05768__I (.I(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05771__I0 (.I(\as2650.regs[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05771__I1 (.I(\as2650.regs[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05772__I (.I(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05773__I (.I(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05775__A2 (.I(\as2650.regs[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05780__A2 (.I(\as2650.regs[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05782__I (.I(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05786__I (.I(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05787__I (.I(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05788__I0 (.I(\as2650.regs[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05788__I1 (.I(\as2650.regs[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05789__I (.I(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05792__I (.I(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05793__I (.I(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05795__A1 (.I(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05797__I (.I(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05801__I (.I(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05803__A2 (.I(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05804__A1 (.I(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05804__A2 (.I(\as2650.regs[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05805__I (.I(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05808__I (.I(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05809__I (.I(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05814__I (.I(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05818__A1 (.I(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05820__I (.I(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05821__I (.I(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05825__I (.I(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05828__I (.I(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05829__I (.I(\as2650.indirect_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05830__A1 (.I(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05830__A2 (.I(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05831__A1 (.I(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05831__A2 (.I(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05831__A3 (.I(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05833__A1 (.I(\as2650.wb_hidden_rom_enable ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05836__I (.I(\as2650.wb_hidden_rom_enable ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05841__A3 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05844__I (.I(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05846__A1 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05847__A1 (.I(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05847__A2 (.I(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05851__I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05856__A1 (.I(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05856__B (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05861__I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05863__B (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05866__I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05867__B (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05872__I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05873__A1 (.I(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05873__B (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05875__A3 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05876__A1 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05879__I (.I(\as2650.extend ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05880__A2 (.I(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05880__A3 (.I(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05880__B (.I(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05881__A3 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05882__A1 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05886__I0 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05886__I1 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05889__A1 (.I(\as2650.indirect_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05889__A2 (.I(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05889__A3 (.I(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05890__A3 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05891__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05895__A1 (.I(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05896__I (.I(\as2650.extend ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05897__A1 (.I(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05897__A2 (.I(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05899__A1 (.I(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05900__A1 (.I(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05900__A2 (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05904__A2 (.I(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05905__A1 (.I(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05908__A2 (.I(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05910__I (.I(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05911__A2 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05912__A1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05912__C (.I(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05913__I (.I(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05915__I (.I(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05919__I (.I(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05920__I (.I(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05921__I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05922__B (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05924__I (.I(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05925__I (.I(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05928__A1 (.I(\as2650.regs[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05929__A2 (.I(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05930__I (.I(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05931__I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05932__B (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05933__C (.I(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05934__I (.I(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05937__A1 (.I(\as2650.regs[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05938__A4 (.I(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05939__I (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05940__A1 (.I(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05940__A2 (.I(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05940__A3 (.I(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05940__A4 (.I(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05942__I (.I(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05943__A1 (.I(\as2650.regs[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05943__A2 (.I(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05943__B2 (.I(\as2650.regs[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05944__A1 (.I(\as2650.regs[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05946__A1 (.I(\as2650.regs[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05947__I (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05950__A1 (.I(\as2650.regs[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05950__B2 (.I(\as2650.regs[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05952__I (.I(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05954__A1 (.I(\as2650.regs[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05957__A1 (.I(\as2650.regs[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05957__A2 (.I(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05960__B (.I(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05961__A4 (.I(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05963__A1 (.I(\as2650.regs[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05963__A2 (.I(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05964__A1 (.I(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05964__A3 (.I(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05967__A1 (.I(\as2650.regs[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05967__A2 (.I(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05972__A1 (.I(\as2650.regs[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05975__A1 (.I(\as2650.regs[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05975__C (.I(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05977__A1 (.I(\as2650.regs[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05978__A1 (.I(\as2650.regs[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05978__A2 (.I(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05983__A1 (.I(\as2650.regs[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05984__A1 (.I(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05988__A1 (.I(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05988__B2 (.I(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05992__A1 (.I(\as2650.regs[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05992__A3 (.I(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05993__A1 (.I(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05995__I (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05997__A1 (.I(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06001__I (.I(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06002__I (.I(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06003__A1 (.I(\as2650.regs[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06004__A1 (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06005__I (.I(\as2650.regs[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06007__A1 (.I(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06007__B2 (.I(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06007__C (.I(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06009__A1 (.I(\as2650.regs[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06010__A1 (.I(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06012__I (.I(\as2650.regs[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06013__A2 (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06015__I (.I(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06016__I (.I(\as2650.regs[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06017__I (.I(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06018__B (.I(\as2650.regs[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06021__I (.I(\as2650.regs[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06025__I (.I(\as2650.regs[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06027__A1 (.I(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06028__I (.I(\as2650.regs[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06031__B1 (.I(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06034__B (.I(\as2650.regs[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06037__I (.I(\as2650.regs[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06038__I (.I(\as2650.regs[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06042__A1 (.I(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06043__I (.I(\as2650.regs[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06048__I (.I(\as2650.regs[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06049__I (.I(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06050__B (.I(\as2650.regs[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06052__I (.I(\as2650.regs[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06053__I (.I(\as2650.regs[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06054__A1 (.I(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06057__A1 (.I(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06060__A1 (.I(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06063__B (.I(\as2650.regs[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06065__I (.I(\as2650.regs[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06066__I (.I(\as2650.regs[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06070__A1 (.I(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06071__I (.I(\as2650.regs[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06075__A4 (.I(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06076__A1 (.I(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06076__A2 (.I(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06077__A1 (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06079__A1 (.I(\as2650.extend ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06081__I (.I(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06082__I (.I(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06084__A1 (.I(\as2650.regs[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06085__A1 (.I(\as2650.regs[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06085__A2 (.I(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06085__C (.I(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06087__A1 (.I(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06089__A4 (.I(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06090__A1 (.I(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06091__A1 (.I(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06093__A1 (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06094__A2 (.I(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06095__A1 (.I(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06096__I (.I(\as2650.indirect_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06097__A1 (.I(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06098__I (.I(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06099__I (.I(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06102__A1 (.I(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06102__A2 (.I(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06106__A1 (.I(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06109__I (.I(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06110__B2 (.I(\as2650.PC[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06111__B2 (.I(\as2650.PC[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06112__A2 (.I(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06112__B1 (.I(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06112__B2 (.I(\as2650.PC[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06114__A2 (.I(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06115__A1 (.I(\as2650.PC[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06115__A2 (.I(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06119__A2 (.I(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06120__A1 (.I(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06120__A2 (.I(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06121__A2 (.I(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06121__B2 (.I(\as2650.PC[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06123__A2 (.I(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06124__I0 (.I(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06124__S (.I(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06127__A2 (.I(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06128__A1 (.I(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06130__A2 (.I(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06130__B1 (.I(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06130__B2 (.I(\as2650.PC[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06133__A2 (.I(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06135__I (.I(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06137__A1 (.I(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06139__A2 (.I(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06141__A1 (.I(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06142__A1 (.I(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06142__A2 (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06146__A4 (.I(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06147__I (.I(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06148__I (.I(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06150__B (.I(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06151__I (.I(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06152__I (.I(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06153__A2 (.I(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06155__A1 (.I(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06156__A1 (.I(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06158__I (.I(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06160__A1 (.I(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06160__A2 (.I(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06162__A2 (.I(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06163__A2 (.I(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06164__A1 (.I(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06168__A1 (.I(\as2650.regs[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06169__A1 (.I(\as2650.regs[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06169__A2 (.I(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06169__B2 (.I(\as2650.regs[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06171__A3 (.I(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06174__A1 (.I(\as2650.regs[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06174__B2 (.I(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06177__A1 (.I(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06177__A2 (.I(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06178__A1 (.I(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06182__A1 (.I(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06183__A2 (.I(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06184__A1 (.I(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06184__A2 (.I(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06186__A1 (.I(\as2650.regs[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06187__A1 (.I(\as2650.regs[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06187__C (.I(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06190__A1 (.I(\as2650.regs[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06192__A1 (.I(\as2650.regs[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06195__A1 (.I(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06197__A1 (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06197__A2 (.I(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06197__B (.I(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06198__A1 (.I(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06201__A1 (.I(\as2650.instruction_args_latch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06202__A1 (.I(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06202__B2 (.I(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06203__A1 (.I(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06205__A1 (.I(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06208__A1 (.I(\as2650.regs[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06208__A2 (.I(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06210__A1 (.I(\as2650.regs[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06210__A2 (.I(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06210__B1 (.I(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06210__B2 (.I(\as2650.regs[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06212__A3 (.I(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06215__A1 (.I(\as2650.regs[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06218__I (.I(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06220__I (.I(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06221__A1 (.I(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06222__A1 (.I(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06223__A2 (.I(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06225__A1 (.I(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06226__I (.I(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06227__A1 (.I(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06228__A2 (.I(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06232__A1 (.I(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06234__A1 (.I(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06235__I (.I(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06239__A2 (.I(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06239__C (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06245__A1 (.I(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06245__A2 (.I(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06247__A1 (.I(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06251__A2 (.I(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06252__A1 (.I(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06253__A1 (.I(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06258__A2 (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06261__A1 (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06265__A1 (.I(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06265__A2 (.I(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06266__A2 (.I(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06268__A1 (.I(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06271__A1 (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06271__A2 (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06272__A1 (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06272__C (.I(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06273__A2 (.I(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06273__C (.I(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06275__S (.I(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06276__A2 (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06280__A1 (.I(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06281__A1 (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06282__A1 (.I(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06284__A1 (.I(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06284__A2 (.I(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__A1 (.I(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06286__A1 (.I(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06289__I (.I(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06291__B2 (.I(\as2650.PC[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06292__A3 (.I(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06296__A1 (.I(\as2650.PC[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06300__A1 (.I(\as2650.indirect_target[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06300__B2 (.I(\as2650.PC[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06301__I (.I(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06302__B2 (.I(\as2650.PC[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06303__B (.I(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06305__A3 (.I(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06307__A1 (.I(\as2650.instruction_args_latch[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06307__A2 (.I(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06310__A1 (.I(\as2650.instruction_args_latch[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06313__A1 (.I(\as2650.instruction_args_latch[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06315__I (.I(\as2650.instruction_args_latch[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06316__I (.I(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06319__A1 (.I(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06320__A3 (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06325__B2 (.I(\as2650.PC[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06327__A1 (.I(\as2650.instruction_args_latch[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06328__A1 (.I(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06330__I (.I(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06332__A1 (.I(\as2650.ivectors_base[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06333__A2 (.I(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06336__A2 (.I(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06336__A3 (.I(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06337__B2 (.I(\as2650.page_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06339__A1 (.I(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06339__A2 (.I(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06340__I (.I(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__A1 (.I(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__A2 (.I(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06342__A1 (.I(\as2650.page_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06343__A1 (.I(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06349__I (.I(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06350__I (.I(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06353__A1 (.I(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06353__A2 (.I(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06354__A1 (.I(\as2650.ivectors_base[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06355__A1 (.I(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06358__I (.I(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06359__A1 (.I(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06360__C (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06361__A3 (.I(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06362__I (.I(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06366__I (.I(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06367__A1 (.I(\as2650.ivectors_base[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06367__A2 (.I(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06368__A1 (.I(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06371__A1 (.I(\as2650.ivectors_base[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06371__A2 (.I(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06372__A2 (.I(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06375__B (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__A2 (.I(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06377__A1 (.I(\as2650.ivectors_base[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06379__A2 (.I(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06381__A1 (.I(\as2650.ivectors_base[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06381__A2 (.I(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06382__A2 (.I(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06385__A1 (.I(\as2650.ivectors_base[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06386__A1 (.I(\as2650.page_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06387__A1 (.I(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06390__B2 (.I(\as2650.page_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06393__A1 (.I(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06394__A1 (.I(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06395__I (.I(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06397__B1 (.I(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06397__B2 (.I(\as2650.page_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06400__I0 (.I(\as2650.instruction_args_latch[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06400__I1 (.I(\as2650.page_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06400__S (.I(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06401__A1 (.I(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06402__A1 (.I(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06403__A1 (.I(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06403__A2 (.I(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06403__A3 (.I(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06404__A1 (.I(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06404__A2 (.I(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06404__B (.I(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06408__A1 (.I(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06408__A2 (.I(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06409__A1 (.I(\as2650.ivectors_base[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06410__A1 (.I(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06417__B (.I(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06418__A2 (.I(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06423__A2 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06424__A1 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06425__I (.I(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06426__I (.I(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06427__I (.I(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06428__A2 (.I(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06430__A2 (.I(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06431__A2 (.I(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06434__A3 (.I(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06439__A2 (.I(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06441__A2 (.I(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06442__A1 (.I(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06443__A2 (.I(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06445__B (.I(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06451__B (.I(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06453__A2 (.I(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06454__A2 (.I(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06455__A2 (.I(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06462__A1 (.I(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06463__A1 (.I(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06466__B (.I(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06467__A1 (.I(\as2650.ivectors_base[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06468__B (.I(_01294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06471__I (.I(\as2650.ivectors_base[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06476__A1 (.I(\as2650.ivectors_base[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06479__B (.I(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06481__A1 (.I(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06485__A1 (.I(\as2650.ivectors_base[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06486__A1 (.I(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06489__A1 (.I(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06489__A2 (.I(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06494__A2 (.I(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06495__I (.I(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06497__I (.I(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06498__I (.I(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06499__I (.I(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06502__I (.I(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06505__I (.I(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06506__I (.I(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06507__I (.I(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06510__I (.I(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06515__I (.I(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06516__I1 (.I(\as2650.regs[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06517__I (.I(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06519__I (.I(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06520__I (.I(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06522__A4 (.I(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06523__I (.I(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06524__I (.I(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06526__I (.I(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06528__A1 (.I(\as2650.warmup[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06528__A2 (.I(\as2650.warmup[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06528__A3 (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06530__I (.I(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06531__I (.I(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06532__I (.I(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06533__I (.I(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06538__I (.I(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06542__I (.I(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06544__I (.I(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06547__A1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06548__A1 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06550__A2 (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06551__A1 (.I(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06551__A2 (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06552__I (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06555__I (.I(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06556__I (.I(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06558__I (.I(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__A1 (.I(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06560__A1 (.I(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06561__A1 (.I(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06562__A2 (.I(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06563__A1 (.I(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06570__I (.I(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06573__A1 (.I(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06573__A2 (.I(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06574__I (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06575__I (.I(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06577__I (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06578__A1 (.I(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06578__A2 (.I(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06578__A3 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06579__I (.I(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06583__A2 (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06585__I (.I(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06587__I (.I(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06588__A2 (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06588__B (.I(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06589__A1 (.I(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06589__A2 (.I(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06590__I (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06592__A1 (.I(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06592__B (.I(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06593__A2 (.I(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06594__A1 (.I(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06594__A2 (.I(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06594__B (.I(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06595__I (.I(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06599__A1 (.I(\as2650.ext_io_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06599__A2 (.I(\as2650.ext_io_addr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06601__A1 (.I(\as2650.io_bus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06602__I (.I(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06603__I (.I(\as2650.ext_io_addr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06604__A1 (.I(\as2650.ext_io_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06606__A1 (.I(\as2650.io_bus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06608__A1 (.I(\as2650.ext_io_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06610__A1 (.I(\as2650.io_bus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06612__A1 (.I(\as2650.warmup[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06612__A2 (.I(\as2650.warmup[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06612__A3 (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06614__I (.I(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06615__I (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06616__I (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06617__I (.I(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06619__I (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06621__I (.I(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06622__A1 (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06622__A4 (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06623__A1 (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06627__I (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06628__I (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06629__I (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06630__A2 (.I(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06630__B2 (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06631__I (.I(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06632__A1 (.I(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06634__I (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06635__I (.I(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06636__I (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06637__A2 (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06637__A3 (.I(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06638__I (.I(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06639__A2 (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06639__A3 (.I(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06640__I (.I(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06644__B (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06645__I (.I(wb_debug_carry));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06649__I (.I(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06651__I (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06652__A1 (.I(wb_debug_cc));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06652__A2 (.I(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06653__A1 (.I(wb_debug_cc));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06653__A2 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06653__B1 (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06653__C (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06654__A1 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06654__A2 (.I(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06658__I (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06660__I (.I(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06661__I (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06662__A1 (.I(wb_debug_cc));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06662__A2 (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06662__B1 (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06662__C (.I(wb_debug_carry));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06663__A1 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06663__A2 (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06665__I (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06667__I (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06670__I (.I(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06671__I (.I(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06672__I (.I(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06674__A2 (.I(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06675__A2 (.I(\as2650.regs[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06676__A2 (.I(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06677__I (.I(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06679__A2 (.I(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06680__A2 (.I(\as2650.regs[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06681__A2 (.I(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06682__A2 (.I(\as2650.regs[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06683__A2 (.I(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06684__A2 (.I(\as2650.regs[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06685__A2 (.I(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06686__I0 (.I(\as2650.regs[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06686__I1 (.I(\as2650.regs[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06686__S (.I(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06688__I0 (.I(\as2650.regs[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06688__I1 (.I(\as2650.regs[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06688__S (.I(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06690__I (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06691__A1 (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06691__A2 (.I(\as2650.regs[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06693__A2 (.I(\as2650.regs[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06695__A2 (.I(\as2650.regs[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06698__I1 (.I(\as2650.regs[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06701__A1 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06701__A2 (.I(\as2650.regs[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06702__A1 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06702__A2 (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06704__A2 (.I(\as2650.regs[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06705__A2 (.I(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__I0 (.I(\as2650.regs[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__I1 (.I(\as2650.regs[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__S (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06708__I0 (.I(\as2650.regs[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06708__I1 (.I(\as2650.regs[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06710__I (.I(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06713__A1 (.I(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06713__A2 (.I(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06714__I (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06716__A2 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06717__A1 (.I(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06718__A1 (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06718__A2 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06719__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06719__A3 (.I(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06720__I (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__A1 (.I(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06723__A2 (.I(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06725__A1 (.I(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06728__I (.I(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06729__A3 (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06733__A1 (.I(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06738__A1 (.I(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06754__I (.I(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06757__B (.I(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06758__A1 (.I(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06759__I (.I(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06762__B (.I(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06763__A1 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06763__A2 (.I(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06764__A1 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06764__A2 (.I(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06764__B (.I(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06765__A2 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06767__A2 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06768__A2 (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06770__A1 (.I(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06772__I (.I(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06774__I (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06777__I (.I(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06778__A1 (.I(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06780__I (.I(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06781__A1 (.I(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06781__A2 (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06782__A2 (.I(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06782__B (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06785__I0 (.I(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06785__I1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06788__I (.I(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06789__A1 (.I(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06790__A1 (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06792__I (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06793__I (.I(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06797__A2 (.I(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06798__A2 (.I(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06798__C (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06799__A1 (.I(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06799__A2 (.I(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06799__B (.I(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06800__A1 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06800__A2 (.I(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06802__A2 (.I(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06803__A1 (.I(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06803__A2 (.I(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06805__A1 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06807__I (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06808__I (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06809__I (.I(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06811__A2 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06812__A2 (.I(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06813__I0 (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06813__S (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__I (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06816__A1 (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06816__A2 (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06819__A1 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06820__I (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06821__I (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06822__I (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06823__A2 (.I(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06824__I (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06825__I0 (.I(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06825__I1 (.I(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06826__A1 (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06828__I (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06830__A1 (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06830__A2 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06833__A1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06841__A1 (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06842__I (.I(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06843__A1 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06844__A1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06845__I (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06847__A2 (.I(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06848__A2 (.I(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06849__A2 (.I(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06851__I (.I(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06854__I (.I(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06856__A1 (.I(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06857__A2 (.I(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06858__A1 (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06859__I (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06860__A1 (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06860__A2 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__A1 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06866__I (.I(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06867__A1 (.I(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06868__A1 (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06869__I (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06871__A2 (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06872__A2 (.I(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06875__A4 (.I(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06876__I (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06878__I (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06880__I (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06881__A1 (.I(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06881__A2 (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06882__I (.I(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06883__A2 (.I(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06884__A1 (.I(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06885__I (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06886__A2 (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06887__A2 (.I(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06889__I (.I(net296));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06891__A1 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06892__I (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06894__I (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06895__A1 (.I(\as2650.instruction_args_latch[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06895__A2 (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06896__A1 (.I(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06897__A1 (.I(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06898__A2 (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06899__A1 (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06900__A1 (.I(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06901__A1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06903__I (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06904__I (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06905__A2 (.I(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06905__A3 (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06906__I (.I(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06907__I (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06908__I (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06909__B (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06910__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06911__I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06912__I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06913__A1 (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06913__A2 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06915__A2 (.I(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06916__A1 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06917__I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06918__A1 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06918__A2 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06921__I (.I(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06922__I (.I(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06923__I0 (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06923__I1 (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06925__I0 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06925__I1 (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06927__I0 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06927__I1 (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06929__I0 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06929__I1 (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06931__I (.I(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06932__I0 (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06932__I1 (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06934__I0 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06934__I1 (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06936__I0 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06936__I1 (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06938__I0 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06938__I1 (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06940__I (.I(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06941__I1 (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06943__I1 (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06945__I0 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06945__I1 (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06947__I0 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06947__I1 (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06949__I (.I(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06950__I1 (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06952__I1 (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06954__I1 (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06956__I1 (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06958__I (.I(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06959__I (.I(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06960__I1 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06962__I1 (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06964__I1 (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06966__I0 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06966__I1 (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06968__I (.I(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06969__I1 (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06971__I0 (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06971__I1 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06973__I0 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06973__I1 (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06975__I0 (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06975__I1 (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06977__I (.I(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06978__I0 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06978__I1 (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06980__I0 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06980__I1 (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06982__I0 (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06982__I1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06984__I0 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06984__I1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06986__I (.I(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06987__I0 (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06987__I1 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06987__S (.I(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06989__I0 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06989__I1 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06989__S (.I(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06991__I0 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06991__I1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06991__S (.I(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06993__I0 (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06993__I1 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06993__S (.I(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06995__I (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06996__I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06997__I (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06998__I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06999__I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07001__A1 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07002__A1 (.I(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07002__A2 (.I(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07003__A3 (.I(net372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07004__I0 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07004__I1 (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07004__S (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07006__I0 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07006__I1 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07006__S (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07008__I0 (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07008__I1 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07008__S (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07010__I (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07011__I (.I(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07013__A1 (.I(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07014__I (.I(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07015__A2 (.I(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07016__I (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07017__I (.I(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07018__A2 (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07019__I (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07020__I (.I(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07021__I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07023__A1 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07023__A2 (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07024__A1 (.I(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07025__A1 (.I(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07025__A2 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07025__B (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07026__A1 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07026__A2 (.I(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__A1 (.I(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07031__A1 (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07031__C (.I(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07033__I (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07034__B (.I(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07035__A2 (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07037__A1 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07037__A2 (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07038__A1 (.I(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07038__A2 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07038__B (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07039__A1 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07039__A2 (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07040__I (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07043__A1 (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07044__A1 (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07044__C (.I(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07045__B (.I(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07046__A2 (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07048__A1 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07048__A2 (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07049__A1 (.I(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07049__A2 (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07049__B (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07050__A1 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07050__A2 (.I(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07052__A1 (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07053__A1 (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07053__C (.I(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07054__B (.I(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07055__I (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07056__I (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07057__I (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07058__I (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07061__I (.I(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07062__A1 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07062__A2 (.I(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07063__I (.I(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07064__A1 (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07067__I (.I(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07068__I (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07069__A1 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07069__A2 (.I(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07070__I (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07071__I (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07072__A1 (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07072__B2 (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07074__A1 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07076__A1 (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07077__I (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07081__A1 (.I(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07081__A2 (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07082__A1 (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07082__B2 (.I(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07084__A1 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07086__I (.I(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07089__A1 (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07092__I (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07093__A2 (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07094__A1 (.I(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07094__B2 (.I(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07098__A1 (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07099__A1 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07099__A2 (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07100__A1 (.I(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07103__I (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07105__I (.I(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07106__I (.I(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07107__A1 (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07108__A1 (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07108__A2 (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07109__I (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07110__A1 (.I(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07114__A1 (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07116__I (.I(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07117__I (.I(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07119__A2 (.I(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07120__A1 (.I(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07123__I (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07126__A1 (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07129__I (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07130__A2 (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07135__A1 (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07137__I (.I(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07138__I (.I(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07140__A2 (.I(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07144__I (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07146__I (.I(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07147__I (.I(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07148__A1 (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07152__I (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07153__A2 (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07154__I (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07159__A1 (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07161__I (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07162__A2 (.I(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07166__I (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07168__A1 (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07170__I (.I(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07171__A2 (.I(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07174__A1 (.I(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07176__A1 (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07177__I (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07178__A2 (.I(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07181__A1 (.I(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07184__A1 (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07184__A2 (.I(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07184__B (.I(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07185__I (.I(\as2650.debug_psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07186__A1 (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07186__A2 (.I(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07187__C (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07188__A2 (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07189__A1 (.I(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07191__I (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07192__I (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07193__I (.I(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07194__A1 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07194__A2 (.I(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07195__A2 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07198__I (.I(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07199__A1 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07199__B (.I(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07200__I (.I(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07201__A1 (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07203__C (.I(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07205__A1 (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07205__B (.I(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07206__I (.I(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07208__I (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07211__A1 (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07211__B (.I(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07216__A1 (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07216__B (.I(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07220__I (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07221__I (.I(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07222__A1 (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07222__B (.I(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07223__I (.I(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07228__A1 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07229__I (.I(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07231__I (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07234__A1 (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07238__A1 (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07242__I (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07243__I (.I(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07244__A1 (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07244__B (.I(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07245__I (.I(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07249__A1 (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07250__I (.I(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07252__I (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07253__B1 (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07255__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07255__B (.I(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07259__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07259__B (.I(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07262__I (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07263__I (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07264__I (.I(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07265__A1 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07265__A2 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07265__B (.I(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07266__I (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07269__I (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07270__A1 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07270__A2 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07270__B (.I(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07271__A1 (.I(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07272__C (.I(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07273__I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__A2 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__B (.I(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07275__A1 (.I(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07276__B1 (.I(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07276__C (.I(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07277__I (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07278__A1 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07278__A2 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07278__B2 (.I(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07279__A1 (.I(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07280__B1 (.I(net392));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07280__C (.I(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07281__A1 (.I(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07281__A2 (.I(net378));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07283__I (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07284__A1 (.I(net334));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07286__I (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07287__A1 (.I(wb_debug_cc));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07288__B (.I(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07289__A1 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07290__A1 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07291__I (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07297__I (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07300__A1 (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07300__A2 (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07303__A1 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07303__A2 (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07305__B (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07306__A1 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07306__A2 (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07306__B (.I(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07307__A1 (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07308__A1 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07308__A2 (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07309__A1 (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07310__B (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07311__I (.I(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07312__A1 (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07312__A2 (.I(net372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07312__B (.I(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07313__A1 (.I(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07313__A2 (.I(net372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07314__A1 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07314__A2 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07314__A3 (.I(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07315__I (.I(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07317__A1 (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07318__A2 (.I(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07318__C (.I(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07320__A1 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07321__A1 (.I(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07321__C (.I(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07325__A1 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07326__A1 (.I(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07326__C (.I(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07327__I (.I(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07328__I (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07329__I (.I(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07331__I (.I(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07332__I (.I(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07333__B (.I(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07338__A1 (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07338__B (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07344__B (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07349__A1 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07349__B (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07351__I (.I(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07353__I (.I(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07354__A1 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07354__B (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07369__I (.I(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07372__I (.I(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07380__B (.I(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07383__B (.I(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07387__B (.I(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07389__I (.I(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07390__I (.I(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07395__I (.I(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07396__B (.I(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07399__I (.I(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07400__I (.I(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07412__I (.I(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07415__I (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07416__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07421__I (.I(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07426__A1 (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07430__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07432__I (.I(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07436__I (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07437__A1 (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07441__I (.I(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07442__A1 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07446__A1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07451__A1 (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07453__I (.I(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07456__I (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07457__A1 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07457__A2 (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07458__A1 (.I(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07461__I (.I(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07462__A1 (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07462__A2 (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07463__A1 (.I(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07467__A1 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07467__A2 (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07468__A1 (.I(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07471__A1 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07471__A2 (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07472__A1 (.I(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07475__A1 (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07475__A2 (.I(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07476__A1 (.I(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07478__A2 (.I(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07479__A1 (.I(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07479__A2 (.I(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07480__A1 (.I(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07482__A1 (.I(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07484__A1 (.I(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07484__B (.I(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07485__A2 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07488__A1 (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07488__A2 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07489__A1 (.I(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__A1 (.I(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__A2 (.I(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07491__I (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07492__I (.I(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07493__A1 (.I(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07493__A2 (.I(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07494__I (.I(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07497__A1 (.I(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07497__A2 (.I(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07498__A1 (.I(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07498__B1 (.I(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07498__B2 (.I(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07499__A1 (.I(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07500__A1 (.I(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07500__A2 (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07501__A1 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07501__A2 (.I(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07504__A1 (.I(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07507__A1 (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07507__A2 (.I(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07509__A1 (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07510__A1 (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07510__A2 (.I(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07512__A1 (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07514__A1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07514__B2 (.I(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07515__A1 (.I(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07516__A1 (.I(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07517__A1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07520__A1 (.I(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07520__A2 (.I(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07521__I (.I(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07522__A1 (.I(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07522__A2 (.I(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07522__B (.I(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07523__A1 (.I(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07527__A2 (.I(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07528__A2 (.I(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07529__A2 (.I(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07531__A2 (.I(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07532__A1 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07532__A3 (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07533__A1 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07534__A1 (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07535__A1 (.I(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07535__A2 (.I(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07536__A2 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07538__I (.I(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07539__I (.I(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__A1 (.I(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__A2 (.I(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__A3 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__A4 (.I(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07542__A1 (.I(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07542__B (.I(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07542__C (.I(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07543__A1 (.I(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07543__A2 (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07545__I (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07547__A1 (.I(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07547__A2 (.I(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07548__A2 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07548__B1 (.I(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07549__I (.I(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07550__A1 (.I(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07551__A1 (.I(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07551__A2 (.I(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07553__I (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07557__I (.I(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07558__A1 (.I(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07558__A2 (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07560__I (.I(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07561__I (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07562__I (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07563__I (.I(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07564__I (.I(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07565__A1 (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07566__A1 (.I(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07566__A2 (.I(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07566__A3 (.I(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07567__I (.I(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07569__I (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07570__A1 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07570__A2 (.I(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07571__I (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07573__I (.I(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07574__I (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07576__A1 (.I(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07577__A1 (.I(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07579__I (.I(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07581__I (.I(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07582__I (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07583__A1 (.I(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07584__I (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07586__I (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07587__I (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07588__I (.I(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07589__I (.I(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07591__A1 (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__A1 (.I(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__A2 (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__A3 (.I(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07594__I (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07596__A1 (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07596__A2 (.I(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07599__A1 (.I(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07600__I (.I(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07601__I1 (.I(\as2650.stack[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07604__I (.I(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07607__A1 (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07609__A1 (.I(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07610__I (.I(\as2650.PC[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07612__I (.I(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07613__I (.I(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07614__I (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07615__I (.I(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07616__I (.I(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07617__A1 (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07620__B (.I(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07621__A2 (.I(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07622__I (.I(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07623__I0 (.I(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07623__I1 (.I(\as2650.stack[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07627__I (.I(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07629__A1 (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07630__A1 (.I(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07631__I (.I(\as2650.PC[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07635__A2 (.I(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07636__B (.I(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07637__A2 (.I(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07638__I (.I(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07639__I1 (.I(\as2650.stack[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07641__A1 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07642__A1 (.I(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07644__I (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07645__I (.I(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07646__A3 (.I(\as2650.PC[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07651__A2 (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07652__I (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07653__I1 (.I(\as2650.stack[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07655__I (.I(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07656__A1 (.I(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07658__A1 (.I(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07659__I (.I(\as2650.PC[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07661__A1 (.I(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07663__A2 (.I(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07665__A1 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07666__I (.I(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07667__I (.I(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07670__I (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07671__A1 (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07672__A1 (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07673__I (.I(\as2650.PC[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07674__I (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07675__I (.I(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07676__A1 (.I(\as2650.PC[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07677__A2 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07678__A1 (.I(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07680__A1 (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07681__I (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07688__A1 (.I(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07689__A1 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07690__I (.I(\as2650.PC[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07692__A1 (.I(\as2650.PC[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07692__A2 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07695__A1 (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07695__A2 (.I(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07696__A1 (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07697__A1 (.I(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07698__I (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07701__I (.I(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07702__A1 (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07703__A1 (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07704__I (.I(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07705__I (.I(\as2650.PC[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07707__A1 (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07707__A3 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07710__I (.I(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07712__I (.I(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07713__A2 (.I(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07714__A1 (.I(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07715__I (.I(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07716__I0 (.I(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07719__A1 (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07721__A1 (.I(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07722__I (.I(\as2650.PC[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07726__I (.I(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07730__C (.I(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07731__A2 (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07732__I (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07733__I (.I(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07734__I0 (.I(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07734__I1 (.I(\as2650.stack[11][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07737__A1 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07738__A1 (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07739__I (.I(\as2650.PC[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07741__A1 (.I(\as2650.PC[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07742__I (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07743__A1 (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07743__A2 (.I(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07744__A1 (.I(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07744__B (.I(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07745__A2 (.I(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07746__I (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07747__I0 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07749__I (.I(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07750__I (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07751__A1 (.I(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07753__I (.I(\as2650.PC[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07755__A2 (.I(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07756__A1 (.I(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07758__A1 (.I(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07759__A2 (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07759__C (.I(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07760__A2 (.I(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07761__I (.I(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07762__I1 (.I(\as2650.stack[11][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07764__I (.I(\as2650.PC[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07766__A1 (.I(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07768__I (.I(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07770__A2 (.I(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07772__I (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07773__A1 (.I(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07775__A2 (.I(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07776__I (.I(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07781__A1 (.I(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07782__A1 (.I(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07783__I (.I(\as2650.PC[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07784__A1 (.I(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07786__A1 (.I(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07788__A1 (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07788__A2 (.I(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__A1 (.I(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__B (.I(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07790__A1 (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07791__I (.I(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07792__I (.I(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07795__I (.I(\as2650.page_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07796__A1 (.I(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07797__I (.I(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07799__A1 (.I(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__A1 (.I(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07801__A2 (.I(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07802__I (.I(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07805__I (.I(\as2650.page_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07806__A1 (.I(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07809__A1 (.I(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07810__A1 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07811__A2 (.I(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07812__I (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07815__I (.I(\as2650.page_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07816__A1 (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07819__A1 (.I(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07820__A1 (.I(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07821__A2 (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07822__I (.I(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07823__I0 (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07826__A1 (.I(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07826__A2 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07827__I (.I(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07829__I (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07830__I (.I(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07832__I (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07833__I (.I(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07834__I (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07835__A2 (.I(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07835__B (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07836__A2 (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07838__I (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07839__I1 (.I(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07841__I0 (.I(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07841__I1 (.I(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07845__I1 (.I(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07847__I (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07848__S (.I(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07850__S (.I(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07852__S (.I(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07854__I0 (.I(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07854__S (.I(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07856__I (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07857__I0 (.I(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07859__I0 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07859__I1 (.I(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07865__I (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07866__S (.I(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07868__S (.I(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07870__S (.I(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07872__I0 (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07872__S (.I(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07875__I (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07876__I1 (.I(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07878__I0 (.I(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07878__I1 (.I(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07882__I1 (.I(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07884__I (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07885__S (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07887__S (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07889__S (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07891__I0 (.I(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07891__S (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07893__I (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07894__I0 (.I(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07896__I0 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07896__I1 (.I(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07902__I (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07903__S (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07905__S (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__S (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07909__I0 (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07909__S (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07916__A1 (.I(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07917__I (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07918__I1 (.I(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07920__I0 (.I(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07926__I (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07927__S (.I(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07929__S (.I(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07931__S (.I(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07933__I0 (.I(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07933__S (.I(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07935__I (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07936__I0 (.I(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07938__I0 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07944__I (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07945__I1 (.I(\as2650.stack[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07945__S (.I(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07947__S (.I(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07949__I1 (.I(\as2650.stack[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07949__S (.I(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07951__I0 (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07951__S (.I(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07953__I (.I(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07956__I (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07957__I0 (.I(\as2650.stack[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07959__I (.I(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07962__I (.I(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07965__I (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07968__I (.I(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07969__I (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__I (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__I0 (.I(\as2650.stack[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07975__I (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07976__I0 (.I(\as2650.stack[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07978__I (.I(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07981__I (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07982__I (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07983__I1 (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07985__I (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07986__I1 (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07988__I (.I(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07989__I1 (.I(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07991__I (.I(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07992__I0 (.I(\as2650.stack[14][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07992__I1 (.I(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07994__I (.I(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07995__I (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07996__S (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07998__I (.I(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__S (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08001__I (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08002__S (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08004__I (.I(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08005__S (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08007__A2 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08008__I (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08010__I (.I(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__I (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08013__I (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__I (.I(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08016__I0 (.I(\as2650.stack[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08016__S (.I(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__S (.I(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08020__S (.I(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08022__I0 (.I(\as2650.stack[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08022__S (.I(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08024__I (.I(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08027__I0 (.I(\as2650.stack[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__I (.I(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08034__I1 (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08036__I1 (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08038__I1 (.I(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08040__I0 (.I(\as2650.stack[13][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08040__I1 (.I(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08042__I (.I(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08043__S (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08045__S (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08047__S (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08049__S (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08051__I (.I(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08052__A1 (.I(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08053__I (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__S (.I(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08056__I (.I(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08057__I1 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08057__S (.I(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08059__I (.I(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08060__I1 (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08060__S (.I(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08062__I (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08063__I1 (.I(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08063__S (.I(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08065__I (.I(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08066__I (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08067__I0 (.I(\as2650.stack[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08069__I (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__I0 (.I(\as2650.stack[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08072__I (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__I0 (.I(\as2650.stack[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08075__I (.I(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08078__I (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__I (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__I1 (.I(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08082__I (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08083__I1 (.I(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__I (.I(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08088__I (.I(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08089__I1 (.I(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08091__I (.I(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08092__I (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08093__S (.I(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08095__I (.I(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08096__I0 (.I(\as2650.stack[12][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08096__S (.I(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08098__I (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08099__S (.I(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08101__I (.I(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08102__S (.I(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08104__I (.I(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08105__A1 (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__I (.I(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08107__S (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__I (.I(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08110__I0 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08110__S (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08112__I (.I(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08113__I0 (.I(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08113__S (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08115__I (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08116__S (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08118__I (.I(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__I (.I(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08122__I (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08125__I (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08128__I (.I(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08131__I (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08132__I (.I(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08133__I0 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08133__S (.I(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__I (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08136__I0 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08136__S (.I(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08138__I (.I(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08139__S (.I(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08141__I (.I(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08142__I0 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08142__S (.I(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08144__I (.I(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08145__I (.I(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08148__I (.I(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08151__I (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__I (.I(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08157__A1 (.I(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08157__A2 (.I(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08158__I (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08159__S (.I(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08161__I0 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08161__S (.I(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08163__I0 (.I(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08163__S (.I(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08165__S (.I(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08167__I (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08170__I1 (.I(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08176__I (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08177__I0 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08179__I0 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08183__I0 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08185__I (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08194__A2 (.I(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08195__I (.I(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__S (.I(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08198__I1 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08198__S (.I(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08200__I1 (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08200__S (.I(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08202__I1 (.I(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08202__S (.I(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08204__I (.I(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08205__I0 (.I(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08207__I0 (.I(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08209__I0 (.I(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08211__I0 (.I(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08213__I (.I(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08214__I1 (.I(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08216__I1 (.I(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08220__I1 (.I(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08222__I (.I(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08223__I0 (.I(\as2650.stack[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08223__S (.I(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08225__I0 (.I(\as2650.stack[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08225__S (.I(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08227__I0 (.I(\as2650.stack[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08227__S (.I(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08229__I0 (.I(\as2650.stack[6][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08229__S (.I(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08232__I (.I(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08233__S (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08235__I1 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08235__S (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08237__I1 (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08237__S (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08239__I1 (.I(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08239__S (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08241__I (.I(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08244__I0 (.I(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08246__I0 (.I(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08250__I (.I(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08251__I1 (.I(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08253__I1 (.I(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08257__I0 (.I(\as2650.stack[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08257__I1 (.I(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08259__I (.I(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08268__A1 (.I(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08269__I (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08270__S (.I(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08272__I0 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08272__S (.I(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08274__I0 (.I(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08274__S (.I(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__S (.I(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08278__I (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08287__I (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08288__I0 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08288__S (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08290__I0 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08290__S (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08292__S (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08294__I0 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08294__S (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08296__I (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08305__A1 (.I(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08306__I (.I(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08307__S (.I(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08309__I1 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08309__S (.I(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08311__I1 (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08311__S (.I(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08313__I1 (.I(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08313__S (.I(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08315__I (.I(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08316__I0 (.I(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08318__I0 (.I(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08320__I0 (.I(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08322__I0 (.I(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08324__I (.I(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08325__I1 (.I(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__I1 (.I(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08331__I0 (.I(\as2650.stack[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08331__I1 (.I(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08333__I (.I(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08340__I0 (.I(\as2650.stack[4][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08343__I (.I(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08344__S (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08346__I0 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08346__S (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08348__I0 (.I(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08348__S (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08350__S (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08352__I (.I(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08355__I1 (.I(\as2650.stack[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08361__I (.I(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08362__I0 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08362__S (.I(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08364__I0 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08364__S (.I(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08366__S (.I(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08368__I0 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08368__S (.I(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08370__I (.I(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08371__S (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08373__S (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08375__S (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08377__S (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08379__I (.I(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08380__I (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08381__I (.I(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08384__I (.I(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08386__I (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08388__A1 (.I(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08388__A2 (.I(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08389__A2 (.I(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08390__A1 (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08390__A2 (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08392__A2 (.I(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08392__A3 (.I(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08393__A1 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08393__A2 (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08395__A1 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08396__A1 (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08396__A2 (.I(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08397__A1 (.I(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08397__A2 (.I(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08398__I (.I(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08399__A2 (.I(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__A2 (.I(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08402__A2 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08402__A3 (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08404__I (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08405__A1 (.I(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08405__A2 (.I(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08405__A3 (.I(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08406__A2 (.I(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08406__A3 (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08407__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08407__A2 (.I(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08408__A2 (.I(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08409__A1 (.I(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08409__A2 (.I(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08409__A3 (.I(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08410__A1 (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08411__A1 (.I(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08412__A1 (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08412__A2 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08412__A3 (.I(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08416__A1 (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08416__A2 (.I(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08417__A1 (.I(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08418__A1 (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08418__A2 (.I(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08418__A4 (.I(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08419__A1 (.I(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08419__A2 (.I(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08420__A1 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08420__A2 (.I(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08420__A3 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08421__A2 (.I(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08422__A1 (.I(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08424__A1 (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08424__A2 (.I(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08427__A3 (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08428__A1 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08428__A2 (.I(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08428__A3 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08429__I (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08431__I (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08432__A1 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08432__A2 (.I(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08437__A3 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08437__A4 (.I(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08438__A2 (.I(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08438__A3 (.I(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08439__A1 (.I(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08440__I (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08441__I (.I(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08446__B2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08449__I (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08450__I (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08451__I (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08452__A1 (.I(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08456__I (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08457__A1 (.I(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08461__I (.I(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08462__I (.I(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08463__A1 (.I(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08463__A2 (.I(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08465__A1 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08465__A2 (.I(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08469__A1 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08473__B (.I(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__A1 (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__I (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08478__A1 (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08478__A2 (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__A1 (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__A3 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08480__A1 (.I(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08480__A2 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08481__A1 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08481__A3 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08486__A1 (.I(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08487__A2 (.I(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__A2 (.I(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08491__A2 (.I(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08492__A2 (.I(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08493__A1 (.I(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08496__A2 (.I(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__A1 (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__A2 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__I (.I(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08500__A1 (.I(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__B (.I(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08502__A1 (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08505__I (.I(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08506__I (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__A1 (.I(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08508__A1 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08509__A1 (.I(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08509__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08510__A1 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08511__B (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08512__A1 (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08512__A2 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__I (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08514__I (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08515__I (.I(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08516__A3 (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__I (.I(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08520__A1 (.I(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08520__A2 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08520__A4 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08521__A1 (.I(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__I (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08525__I (.I(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__A1 (.I(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__B (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__C (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08527__I (.I(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08528__A1 (.I(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08528__B1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08528__B2 (.I(\as2650.regs[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08529__A2 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08531__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08531__B2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__A1 (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08534__A1 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08535__I (.I(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08536__I (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08537__A2 (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08538__A1 (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08538__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08539__I (.I(_02979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08540__A1 (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08540__A2 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08541__I (.I(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08542__I (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__A1 (.I(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__A2 (.I(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08544__B (.I(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08545__A1 (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08545__A2 (.I(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08546__B (.I(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__A1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08550__A2 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08557__A2 (.I(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08560__A1 (.I(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08562__A1 (.I(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08562__C (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08563__A1 (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__A1 (.I(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08566__I (.I(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08569__I (.I(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08570__A2 (.I(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08574__A1 (.I(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08574__A2 (.I(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08576__A2 (.I(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08577__A1 (.I(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08578__A1 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08580__A2 (.I(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08581__A1 (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08581__A2 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08583__C (.I(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08584__A1 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08585__A1 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08586__A1 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08586__A2 (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08588__A1 (.I(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08590__A1 (.I(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__I (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08592__A1 (.I(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08593__A1 (.I(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08594__I (.I(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08595__I (.I(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__I (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08597__I (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08598__A1 (.I(\as2650.regs[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08598__B1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08599__A2 (.I(_03035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08600__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08600__C1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08601__A1 (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08601__A2 (.I(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08602__I (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08603__A2 (.I(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08604__I (.I(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08608__I (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08610__A1 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08611__A2 (.I(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08612__I0 (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08612__I1 (.I(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08612__S (.I(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08618__I0 (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08618__I1 (.I(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08618__S (.I(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__A1 (.I(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08625__A1 (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08626__B (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08627__A1 (.I(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08629__I (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08631__I (.I(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__A1 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08634__A1 (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08636__A1 (.I(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08638__A1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08640__A1 (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08641__A2 (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08643__B (.I(_02979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08644__I (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08645__A1 (.I(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08646__A1 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08647__I (.I(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08648__I (.I(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__I (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08650__A1 (.I(\as2650.regs[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08650__B1 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08651__A2 (.I(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08652__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08652__C1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08653__I0 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08653__I1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__I (.I(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__A1 (.I(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08657__A2 (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08659__A1 (.I(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08659__A2 (.I(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08660__A2 (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08665__A1 (.I(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08665__A2 (.I(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__A1 (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08672__A1 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08673__A1 (.I(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__A1 (.I(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__A1 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__A2 (.I(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__B (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__A1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08682__A1 (.I(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__A1 (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__A1 (.I(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08688__A1 (.I(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__A1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08690__A1 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08691__A1 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08691__A2 (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08693__A1 (.I(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__I (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__A1 (.I(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08697__I0 (.I(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08698__I (.I(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08699__I (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__I (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08701__A1 (.I(\as2650.regs[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08701__B1 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08702__A2 (.I(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08703__I (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08705__B2 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08707__I (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08709__I0 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08710__A1 (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08710__C (.I(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08711__A1 (.I(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08712__A1 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08715__A1 (.I(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08716__A2 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08717__A1 (.I(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08718__A2 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08723__A1 (.I(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__I (.I(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08733__A1 (.I(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08734__B (.I(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08735__A1 (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08739__A2 (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08741__I0 (.I(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08741__S (.I(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08743__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08744__I (.I(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08745__A1 (.I(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08745__A2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08748__A2 (.I(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08749__I (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08750__I (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08751__I (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08752__B1 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08753__A2 (.I(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08755__B2 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08758__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__I (.I(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08760__I (.I(_02979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08761__I0 (.I(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08761__I1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__I0 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__I1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__S (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__A1 (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08775__A1 (.I(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08776__A1 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08780__I (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08783__A1 (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08784__A1 (.I(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08786__C (.I(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08787__A1 (.I(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08788__A1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08789__A2 (.I(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08793__A1 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08793__C (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08794__A2 (.I(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__I (.I(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__I (.I(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__I (.I(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08798__A2 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08798__B1 (.I(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08799__A2 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08803__A1 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__I (.I(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08805__I (.I(_03240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08808__A1 (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08808__A2 (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08809__A1 (.I(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08809__A2 (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08811__A2 (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__A1 (.I(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__A2 (.I(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08821__A1 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__A1 (.I(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08827__A1 (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08827__B2 (.I(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08828__A1 (.I(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08829__A1 (.I(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08829__A2 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08831__A1 (.I(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08832__A2 (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__A1 (.I(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__A1 (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__A1 (.I(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08838__A1 (.I(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08841__A1 (.I(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08842__A1 (.I(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08842__C (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08844__A1 (.I(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08846__A1 (.I(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08846__C (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08847__A2 (.I(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08848__I (.I(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__I (.I(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__I (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08851__A1 (.I(\as2650.regs[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08851__A2 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08851__B1 (.I(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08856__I (.I(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__A2 (.I(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08858__A1 (.I(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__I0 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__I1 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__I0 (.I(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__I1 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__S (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__A1 (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__B2 (.I(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08873__A1 (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08875__A1 (.I(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08877__A2 (.I(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08878__A2 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08878__B (.I(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__A1 (.I(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__A1 (.I(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__A1 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08887__A2 (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08890__A1 (.I(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08891__A2 (.I(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08892__I (.I(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08893__I (.I(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08894__I (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08895__I (.I(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08896__A1 (.I(\as2650.regs[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08896__A2 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08896__B1 (.I(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08899__I (.I(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__I1 (.I(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__S (.I(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08902__S (.I(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08904__S (.I(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08906__S (.I(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08908__I (.I(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08909__I1 (.I(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08909__S (.I(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__I1 (.I(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__S (.I(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08913__I1 (.I(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08913__S (.I(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08915__I1 (.I(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08915__S (.I(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08917__I (.I(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08918__I0 (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08920__I0 (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08922__I0 (.I(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08924__I0 (.I(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08926__I (.I(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08927__S (.I(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08929__I1 (.I(\as2650.stack[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08929__S (.I(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08931__S (.I(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08933__I1 (.I(\as2650.stack[1][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08933__S (.I(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08935__I (.I(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08937__B (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08938__A1 (.I(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08938__A2 (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08940__A1 (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08941__I (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__A2 (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08946__A1 (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08949__B (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08951__A1 (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08954__B (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08955__I (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08957__A1 (.I(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08960__I (.I(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08961__I (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08962__I (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08965__I (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08966__A1 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08967__I (.I(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08968__I (.I(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08970__A1 (.I(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08971__I (.I(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08972__A1 (.I(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08974__A1 (.I(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08974__A3 (.I(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08974__B (.I(\as2650.instruction_args_latch[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08975__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08977__A1 (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08977__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__A1 (.I(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__A2 (.I(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__A3 (.I(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__B1 (.I(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__I (.I(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__A1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__B1 (.I(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08982__A1 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08982__A2 (.I(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08983__I (.I(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__A2 (.I(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08986__A2 (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08988__I (.I(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08990__A1 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08990__A2 (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08990__A3 (.I(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08991__A2 (.I(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08992__B1 (.I(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08993__B (.I(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08995__A1 (.I(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__B (.I(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08997__A1 (.I(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08997__A3 (.I(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08997__B (.I(\as2650.instruction_args_latch[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08998__A2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08999__A1 (.I(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08999__A3 (.I(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09001__I (.I(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09002__A3 (.I(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09003__I (.I(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__A1 (.I(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__A2 (.I(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__A3 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__A4 (.I(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09006__I (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09007__A1 (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09008__A1 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09009__I (.I(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09010__A1 (.I(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09011__A2 (.I(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09011__B2 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09012__A1 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09012__A2 (.I(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09012__B (.I(\as2650.instruction_args_latch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09013__A2 (.I(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09013__A3 (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09013__A4 (.I(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09015__I (.I(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__B2 (.I(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09017__B (.I(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09019__I (.I(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09020__I0 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09020__I1 (.I(\as2650.instruction_args_latch[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09020__S (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09025__A1 (.I(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09025__A2 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09026__I (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09027__I0 (.I(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09027__S (.I(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09028__A1 (.I(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09028__B1 (.I(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09029__B2 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09030__I0 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09031__B2 (.I(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09032__B (.I(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__I (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09035__I (.I(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09036__I (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09037__I (.I(\as2650.instruction_args_latch[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09038__A1 (.I(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09039__A1 (.I(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09043__A1 (.I(_03448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09046__A1 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09047__I (.I(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09049__I (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09051__A1 (.I(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09052__A1 (.I(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09054__B2 (.I(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09056__A1 (.I(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09057__I (.I(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09059__B (.I(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09062__I (.I(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09063__I (.I(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09064__I (.I(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09066__I (.I(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09067__A1 (.I(\as2650.instruction_args_latch[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09068__A1 (.I(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09069__A1 (.I(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__A1 (.I(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__A2 (.I(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__A3 (.I(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__B1 (.I(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__B2 (.I(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09076__A2 (.I(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09077__A1 (.I(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09079__B (.I(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__A1 (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__A2 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09083__A1 (.I(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09084__A1 (.I(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09087__A2 (.I(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09089__A2 (.I(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09089__A3 (.I(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09090__A2 (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09091__A1 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09092__A1 (.I(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09092__A2 (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09093__B1 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09093__B2 (.I(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09094__A2 (.I(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09095__A1 (.I(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__B (.I(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09099__I (.I(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__A1 (.I(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09102__A2 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09103__A2 (.I(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__A2 (.I(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09105__A2 (.I(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09107__A1 (.I(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09108__A1 (.I(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09108__A2 (.I(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09108__B (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09109__B2 (.I(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09110__A2 (.I(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09111__A1 (.I(_03240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09111__A2 (.I(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09113__B (.I(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09115__I (.I(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09116__I (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09120__A2 (.I(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09123__A1 (.I(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09123__A2 (.I(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09123__B (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09126__A1 (.I(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09126__A2 (.I(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__B2 (.I(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09128__B (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__A1 (.I(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09133__I (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09138__A1 (.I(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09138__A2 (.I(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09138__B (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09140__I (.I(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09141__A1 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09141__A2 (.I(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09141__B2 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__A2 (.I(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__B (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09143__I (.I(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09144__I (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09145__I (.I(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09147__I (.I(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09148__I (.I(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09149__A1 (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09149__A2 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09150__A1 (.I(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09153__I (.I(net296));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09154__A2 (.I(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09156__B1 (.I(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09157__A1 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09158__B2 (.I(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09160__I (.I(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__A1 (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09166__A1 (.I(\as2650.indirect_target[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09167__A2 (.I(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09167__A3 (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09168__I (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09169__A1 (.I(\as2650.indirect_target[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09169__B1 (.I(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09169__B2 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09171__A1 (.I(\as2650.instruction_args_latch[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09172__A1 (.I(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09176__A1 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09177__A1 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09180__B2 (.I(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09181__A1 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09185__A1 (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09187__A1 (.I(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09187__A2 (.I(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09188__B2 (.I(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09189__A1 (.I(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09190__B2 (.I(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09192__I (.I(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09193__A2 (.I(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09193__B2 (.I(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09194__I (.I(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09195__I (.I(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09196__A1 (.I(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09197__A1 (.I(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09197__A2 (.I(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09197__B (.I(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09199__A1 (.I(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09201__I (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09202__I (.I(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09203__I0 (.I(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09203__I1 (.I(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09203__S (.I(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09204__B2 (.I(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09205__A1 (.I(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09206__A1 (.I(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09207__A1 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09208__A1 (.I(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09208__B (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09209__A2 (.I(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09209__A3 (.I(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09210__I (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09211__B (.I(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09213__I (.I(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09214__A1 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09214__A2 (.I(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09215__A2 (.I(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09216__A1 (.I(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09216__A2 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09217__I (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09218__A2 (.I(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09220__A2 (.I(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09221__A1 (.I(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__B1 (.I(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09226__A1 (.I(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09227__A1 (.I(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09227__A2 (.I(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09227__B1 (.I(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09228__A1 (.I(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09229__I (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09230__I (.I(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09231__A1 (.I(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09231__A2 (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09232__I (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09233__A1 (.I(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09233__A2 (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09234__A1 (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09236__A1 (.I(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09236__A3 (.I(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09237__B (.I(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09238__A1 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09238__B (.I(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09239__B (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09240__I (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09241__I (.I(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09242__I (.I(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09244__I (.I(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09245__A1 (.I(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09246__A2 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09247__A1 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09247__A2 (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09248__A3 (.I(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09249__A1 (.I(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09249__A3 (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09251__I (.I(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09253__A1 (.I(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09253__A2 (.I(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09253__B (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09254__I (.I(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09255__I (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09256__I (.I(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09257__A1 (.I(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09257__A3 (.I(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09258__A1 (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09260__I (.I(\as2650.warmup[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09261__A1 (.I(\as2650.warmup[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09261__B (.I(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09262__A1 (.I(\as2650.warmup[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09262__A2 (.I(\as2650.warmup[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09263__A1 (.I(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09265__I (.I(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09267__A1 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09267__A2 (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09269__A1 (.I(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09270__A1 (.I(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09271__I (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09273__I (.I(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09274__A1 (.I(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09274__B2 (.I(\as2650.instruction_args_latch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09276__I (.I(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09277__A1 (.I(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09279__A1 (.I(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09281__I (.I(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09282__I (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09284__A1 (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09286__A2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09287__I (.I(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09288__I (.I(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09289__A1 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09291__I (.I(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09292__I (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09293__A1 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__A2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09296__I (.I(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09297__A1 (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09300__I (.I(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09301__I (.I(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09302__A1 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09302__A2 (.I(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09303__A1 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09303__A2 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09303__A3 (.I(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09304__I (.I(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09305__A1 (.I(\as2650.instruction_args_latch[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09306__I (.I(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09307__A1 (.I(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09308__B (.I(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09309__A1 (.I(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09309__B2 (.I(\as2650.instruction_args_latch[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09310__A1 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09311__A1 (.I(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09311__B2 (.I(\as2650.instruction_args_latch[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09312__A1 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09313__A1 (.I(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09313__B2 (.I(\as2650.instruction_args_latch[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09314__A1 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09315__I (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09316__I (.I(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09317__I (.I(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09318__A1 (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09318__B2 (.I(\as2650.instruction_args_latch[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09320__A1 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09320__B2 (.I(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09322__A1 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09324__A1 (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09324__B2 (.I(\as2650.instruction_args_latch[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09326__I (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09327__I (.I(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09328__B (.I(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09329__I (.I(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09331__I (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09333__A1 (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09333__B (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09335__A2 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09335__A3 (.I(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09335__B2 (.I(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09337__B (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09337__C (.I(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09342__A1 (.I(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09342__A2 (.I(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09343__A1 (.I(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09343__A2 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09343__B (.I(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09345__A2 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09348__A1 (.I(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09348__A2 (.I(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09349__A4 (.I(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09353__I (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09354__A1 (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09354__B (.I(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09356__A1 (.I(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09356__A2 (.I(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09356__A3 (.I(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09357__A2 (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09357__B1 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09357__C2 (.I(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09358__A2 (.I(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09360__I (.I(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__A1 (.I(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__A2 (.I(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__C (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09364__A2 (.I(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09365__A1 (.I(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09366__A2 (.I(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09369__A1 (.I(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09371__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09372__I (.I(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09373__A1 (.I(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09373__A2 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09373__A3 (.I(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09374__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09375__A1 (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09375__A2 (.I(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09376__A1 (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09376__A3 (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09376__A4 (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09377__I (.I(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09378__A1 (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09378__A2 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09379__I (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09381__A2 (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09381__B (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09381__C (.I(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09382__A1 (.I(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09383__B (.I(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09384__A1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09385__I (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09386__I (.I(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09387__I (.I(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09388__I (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09389__A2 (.I(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09390__I (.I(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09391__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09391__C (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09392__I (.I(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09393__A2 (.I(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09394__I (.I(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09395__A1 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09395__C (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09396__I (.I(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09397__A2 (.I(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09398__A1 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09398__C (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09399__I (.I(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09400__I (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09401__A2 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09402__A1 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09402__C (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09403__I (.I(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09404__I (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09405__A2 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09406__A1 (.I(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09406__C (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09407__I (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09408__A2 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09409__I (.I(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09410__A1 (.I(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09410__C (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09411__I (.I(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09412__A2 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09413__A1 (.I(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09413__C (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09415__A2 (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__C (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09417__I (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09420__I (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09421__I (.I(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09422__A1 (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09425__A1 (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09426__A1 (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09426__A2 (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09428__A1 (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09429__A1 (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09429__A2 (.I(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09431__A1 (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09431__A2 (.I(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09432__A1 (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09432__A2 (.I(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09434__A1 (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09434__A2 (.I(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09435__A2 (.I(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09435__C (.I(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09438__A1 (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09438__A2 (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09440__A1 (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09440__A2 (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09442__A1 (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09444__A1 (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09446__A1 (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09449__A1 (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09451__A1 (.I(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09451__A2 (.I(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09452__A2 (.I(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09453__A2 (.I(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09455__A1 (.I(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09455__A2 (.I(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09457__B (.I(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09460__A1 (.I(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09460__A2 (.I(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09461__A1 (.I(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09461__A2 (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09462__I (.I(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09463__A1 (.I(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09465__I (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09466__I (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09467__I (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09468__I (.I(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09470__A1 (.I(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09470__A2 (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09471__I (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09472__I (.I(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09473__I (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09474__I (.I(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09475__I (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09477__I (.I(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09478__I (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09484__A3 (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09485__A2 (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09486__I (.I(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09487__I (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09488__I (.I(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09489__I (.I(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09492__B2 (.I(\as2650.stack[12][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09493__I (.I(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09498__I (.I(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09502__A1 (.I(\as2650.stack[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09502__A2 (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09502__B1 (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__B (.I(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09505__A2 (.I(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09505__B1 (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__A1 (.I(\as2650.stack[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__A2 (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__B1 (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09507__A1 (.I(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09511__A1 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09511__A2 (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09512__A1 (.I(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09512__A2 (.I(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09512__C (.I(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09513__A2 (.I(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09514__A1 (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09516__A1 (.I(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09516__A2 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09518__I (.I(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09520__I (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09521__A1 (.I(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09522__I (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__A1 (.I(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__A2 (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09524__A1 (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09526__B2 (.I(\as2650.stack[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09529__A1 (.I(\as2650.stack[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09530__A1 (.I(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09534__A3 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09537__A1 (.I(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09538__A1 (.I(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__I0 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__I1 (.I(\as2650.page_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__A1 (.I(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__B2 (.I(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09542__I (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09543__A1 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09543__B (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__A1 (.I(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__A2 (.I(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__C (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__A2 (.I(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09547__I1 (.I(\as2650.page_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09547__S (.I(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09549__A2 (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09549__B1 (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09550__A1 (.I(\as2650.stack[1][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09550__A2 (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09550__B1 (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09551__A1 (.I(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09552__A2 (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09552__B1 (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09552__B2 (.I(\as2650.stack[4][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__A1 (.I(\as2650.stack[6][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__A2 (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09558__A1 (.I(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__I0 (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__I1 (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09565__A1 (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09565__B2 (.I(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__A1 (.I(\as2650.instruction_args_latch[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__A2 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__B (.I(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09572__B (.I(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09573__A1 (.I(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09575__A1 (.I(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__A1 (.I(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09583__A2 (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09583__B (.I(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09588__A2 (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09588__B (.I(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09589__I (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09590__I (.I(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09591__A2 (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09591__A4 (.I(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__A1 (.I(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__A2 (.I(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09596__A1 (.I(\as2650.ivectors_base[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09597__I (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09598__I (.I(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09599__A1 (.I(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09600__A1 (.I(\as2650.ivectors_base[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09601__A1 (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09602__A1 (.I(\as2650.ivectors_base[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09603__A1 (.I(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09604__A1 (.I(\as2650.ivectors_base[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09605__A1 (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__A1 (.I(\as2650.ivectors_base[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09609__I (.I(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09610__A1 (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09611__A1 (.I(\as2650.ivectors_base[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09612__A1 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__A1 (.I(\as2650.ivectors_base[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09614__A1 (.I(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09615__A1 (.I(\as2650.ivectors_base[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09616__A1 (.I(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09619__A1 (.I(\as2650.ivectors_base[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09620__I (.I(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09621__A1 (.I(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09622__A1 (.I(\as2650.ivectors_base[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09623__A1 (.I(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09624__A1 (.I(\as2650.ivectors_base[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__A1 (.I(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09626__A1 (.I(\as2650.ivectors_base[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09627__A1 (.I(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09629__I (.I(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09630__I (.I(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__A1 (.I(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__A2 (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09632__I (.I(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09633__A2 (.I(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09633__B (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__A1 (.I(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09635__I (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__I (.I(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09638__I (.I(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09639__A1 (.I(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09639__A2 (.I(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__A1 (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09641__I (.I(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09642__I (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09643__A2 (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09643__B1 (.I(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09643__B2 (.I(\as2650.stack[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09646__B1 (.I(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__A1 (.I(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09648__I (.I(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__A1 (.I(\as2650.stack[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__B1 (.I(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09650__A1 (.I(\as2650.stack[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09650__A2 (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09650__B1 (.I(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09653__I (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09656__I (.I(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09657__I (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09658__A2 (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09658__B1 (.I(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09660__A2 (.I(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09660__B1 (.I(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__A1 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__B (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09662__I (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__I (.I(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09664__I (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09665__I (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09666__I (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09668__A1 (.I(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09668__A2 (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09668__B1 (.I(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09668__B2 (.I(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__I (.I(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09672__I (.I(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__A1 (.I(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__A2 (.I(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__B1 (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__B2 (.I(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09674__A1 (.I(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09676__A1 (.I(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09676__A2 (.I(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09677__A1 (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09678__I (.I(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09679__C (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09680__A1 (.I(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09680__A2 (.I(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09681__A1 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09682__I (.I(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09683__I (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09684__A1 (.I(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09685__A1 (.I(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09685__B (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09686__I (.I(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09687__A1 (.I(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09689__I (.I(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09692__A1 (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09693__A2 (.I(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09694__B2 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09695__A1 (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__I (.I(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09697__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09697__A2 (.I(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09697__C (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__A1 (.I(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09701__A1 (.I(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09701__B (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09702__A1 (.I(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09702__A2 (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09702__A3 (.I(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09703__A2 (.I(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09705__A1 (.I(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09705__A2 (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09708__I (.I(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__A1 (.I(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__A2 (.I(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__B1 (.I(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__B2 (.I(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09714__I (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09715__I (.I(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09716__A2 (.I(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09716__B1 (.I(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09717__A1 (.I(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09719__I (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09720__I (.I(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09721__A2 (.I(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09721__B1 (.I(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09724__A2 (.I(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09724__B1 (.I(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09725__A1 (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09727__I (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09730__A2 (.I(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09730__B1 (.I(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09730__B2 (.I(\as2650.stack[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09731__I (.I(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09732__I (.I(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09734__A1 (.I(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09736__A2 (.I(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09736__B1 (.I(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09737__A1 (.I(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09738__A1 (.I(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09739__A1 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__A1 (.I(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__A2 (.I(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__C (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09744__A2 (.I(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09745__A1 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09747__A1 (.I(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09749__A2 (.I(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09750__A1 (.I(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09751__A1 (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09752__A1 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09753__A1 (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09754__A1 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09754__A2 (.I(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09754__C (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09755__I (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09756__I (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09757__A1 (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09760__I (.I(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09761__I (.I(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09763__I (.I(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09765__A2 (.I(_03448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09766__I (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09769__I (.I(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09770__I (.I(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09771__B2 (.I(\as2650.stack[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09773__I (.I(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09775__A1 (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09779__A1 (.I(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09781__I (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09783__I (.I(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09785__I (.I(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09786__I (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09787__I (.I(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09788__A2 (.I(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09788__B1 (.I(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09790__A2 (.I(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09790__B1 (.I(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09791__A1 (.I(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09791__B (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09792__I (.I(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09793__I (.I(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09794__I (.I(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09795__A2 (.I(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09795__B1 (.I(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09796__I (.I(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09797__I (.I(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09798__A2 (.I(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09798__B1 (.I(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09799__A1 (.I(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09800__A1 (.I(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09800__B1 (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09802__A1 (.I(_03448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09802__A2 (.I(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09803__A1 (.I(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09803__A2 (.I(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09805__I (.I(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09806__A2 (.I(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09808__A1 (.I(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09809__A1 (.I(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__A1 (.I(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09811__A2 (.I(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09813__I (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09814__A1 (.I(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09815__I (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09816__I (.I(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__A1 (.I(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__A2 (.I(_03448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09818__I (.I(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09820__B (.I(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09821__I (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09822__A1 (.I(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09824__A1 (.I(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09826__I (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09827__A1 (.I(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09827__B (.I(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09829__I (.I(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09832__I (.I(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09833__I (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09836__I (.I(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09840__A1 (.I(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09841__I (.I(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09842__A1 (.I(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09842__A2 (.I(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09842__B1 (.I(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09842__B2 (.I(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09843__A2 (.I(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09843__B1 (.I(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09844__A1 (.I(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09845__A2 (.I(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09845__B1 (.I(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__A2 (.I(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__B1 (.I(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09847__A1 (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09849__A2 (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09849__B1 (.I(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09849__B2 (.I(\as2650.stack[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09851__A1 (.I(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__A1 (.I(\as2650.stack[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09853__A2 (.I(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09853__B1 (.I(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09854__A1 (.I(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09855__A1 (.I(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09856__A1 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09857__A2 (.I(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09858__I (.I(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09860__A1 (.I(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09861__A1 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09862__A2 (.I(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09863__A1 (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09864__I (.I(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09865__A1 (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09865__C (.I(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09866__A2 (.I(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09867__A1 (.I(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09868__A1 (.I(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__A1 (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09870__A2 (.I(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09871__A1 (.I(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09872__A2 (.I(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09872__B (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09873__B (.I(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09876__A1 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09876__A2 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09876__C (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09877__A1 (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09881__I (.I(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09882__A2 (.I(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09882__B1 (.I(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09883__I (.I(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09884__I (.I(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09885__A1 (.I(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09887__B2 (.I(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09888__I (.I(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09889__I (.I(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09890__A1 (.I(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09890__A2 (.I(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09890__B1 (.I(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09891__A1 (.I(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09893__A2 (.I(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09893__B1 (.I(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09896__B2 (.I(\as2650.stack[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09897__A2 (.I(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09897__B1 (.I(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09898__A1 (.I(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09900__S (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09901__A2 (.I(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09903__A1 (.I(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09903__A2 (.I(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09905__I (.I(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09906__A1 (.I(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09907__A1 (.I(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09907__A2 (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09909__A2 (.I(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09910__A1 (.I(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09911__A1 (.I(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09912__S (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09913__I (.I(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__A1 (.I(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__B (.I(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09916__I (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09917__A1 (.I(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09917__C (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09919__A1 (.I(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09920__A1 (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09920__B (.I(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09924__A2 (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09926__A2 (.I(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09927__I (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09928__A2 (.I(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09928__B1 (.I(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09929__A1 (.I(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09929__A2 (.I(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09929__B1 (.I(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__A1 (.I(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09931__A1 (.I(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09931__A2 (.I(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09931__B1 (.I(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09931__B2 (.I(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09932__A1 (.I(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09932__A2 (.I(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09932__B1 (.I(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09932__B2 (.I(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09933__A1 (.I(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09935__A2 (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09935__B1 (.I(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09936__A1 (.I(\as2650.stack[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09936__A2 (.I(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09936__B1 (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09937__A1 (.I(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09938__A1 (.I(\as2650.stack[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09938__A2 (.I(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09938__B1 (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09938__B2 (.I(\as2650.stack[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09939__A1 (.I(\as2650.stack[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09939__A2 (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09939__B1 (.I(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09939__B2 (.I(\as2650.stack[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09940__A1 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09941__A1 (.I(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09942__A1 (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09943__A2 (.I(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09945__A1 (.I(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__A1 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09947__A2 (.I(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09949__A1 (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09949__B (.I(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09949__C (.I(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__A2 (.I(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09951__A1 (.I(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09952__I (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09953__A1 (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09954__A1 (.I(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09955__B (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09957__A1 (.I(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09957__A2 (.I(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09957__B (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09959__A1 (.I(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09959__A2 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09959__C (.I(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09960__I (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09962__A1 (.I(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09962__A2 (.I(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09962__B1 (.I(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09963__A1 (.I(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09964__A1 (.I(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09964__A2 (.I(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09964__B1 (.I(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09964__B2 (.I(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09965__A1 (.I(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09965__A2 (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09966__A1 (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09968__A2 (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09969__A1 (.I(\as2650.stack[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09969__A2 (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09969__B1 (.I(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09970__A1 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__A2 (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__B1 (.I(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__B2 (.I(\as2650.stack[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09972__A1 (.I(\as2650.stack[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09972__A2 (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09973__A1 (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09974__A1 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09975__A1 (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09976__A1 (.I(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09976__A2 (.I(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09977__A1 (.I(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09978__A1 (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09978__A2 (.I(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09980__A1 (.I(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09980__A2 (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09981__A1 (.I(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09982__A1 (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09982__A2 (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09983__A2 (.I(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__A1 (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__C (.I(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09985__A1 (.I(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09986__A1 (.I(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09986__A2 (.I(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09986__B (.I(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09988__B (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09989__I (.I(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09990__A1 (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09991__A1 (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09994__A1 (.I(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09994__B2 (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09994__C (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09995__A1 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09995__A2 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09996__A2 (.I(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09997__A1 (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09997__A2 (.I(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09999__A1 (.I(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10000__A1 (.I(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__I (.I(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10003__A2 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10003__B1 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10004__A2 (.I(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10004__B1 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10005__A1 (.I(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10006__A2 (.I(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10006__B1 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10007__A2 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10007__B1 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10008__A1 (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10008__A2 (.I(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10010__I (.I(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10011__I (.I(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10014__A2 (.I(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10014__B1 (.I(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10014__B2 (.I(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10016__A1 (.I(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10016__A2 (.I(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10016__B1 (.I(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10017__A1 (.I(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10017__B (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10018__A2 (.I(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10018__B1 (.I(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10019__A1 (.I(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10019__A2 (.I(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10019__B1 (.I(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10020__A1 (.I(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10021__A1 (.I(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10022__A1 (.I(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10022__A2 (.I(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10023__A1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10023__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10024__A1 (.I(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10025__A1 (.I(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10026__A2 (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10027__A1 (.I(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10027__A2 (.I(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10028__A1 (.I(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10028__C (.I(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__A1 (.I(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__A2 (.I(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__B (.I(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10030__A1 (.I(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10031__B (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10032__A1 (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10033__A1 (.I(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10034__B (.I(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10036__B1 (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10036__B2 (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10037__A2 (.I(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10038__A1 (.I(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10039__B (.I(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10041__A3 (.I(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10044__A1 (.I(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10045__B2 (.I(\as2650.stack[11][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10047__A1 (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10051__A1 (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10053__A2 (.I(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10053__B1 (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10055__A2 (.I(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10055__B1 (.I(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__A1 (.I(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__B (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10057__A2 (.I(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10057__B1 (.I(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10058__A2 (.I(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10058__B1 (.I(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10059__A1 (.I(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10060__A1 (.I(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10060__B1 (.I(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10061__A1 (.I(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10061__A2 (.I(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10062__A1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10062__A2 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10063__A1 (.I(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10064__A1 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10065__A2 (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10067__A1 (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10067__C (.I(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10068__A1 (.I(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10068__A2 (.I(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10068__B (.I(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10070__B (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__A1 (.I(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__A2 (.I(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10072__A1 (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10072__C (.I(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10073__A1 (.I(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10074__I (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10075__A1 (.I(\as2650.instruction_args_latch[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10075__B (.I(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10077__A1 (.I(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10078__A1 (.I(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10079__A1 (.I(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10080__B (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10081__A2 (.I(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10081__B (.I(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10083__A2 (.I(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10085__A1 (.I(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10087__A2 (.I(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10087__B1 (.I(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10088__A2 (.I(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10088__B1 (.I(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10089__A1 (.I(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10090__A2 (.I(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10090__B1 (.I(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10091__A2 (.I(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10091__B1 (.I(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10092__A1 (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10093__A1 (.I(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10094__A2 (.I(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10094__B1 (.I(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__A2 (.I(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__B1 (.I(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10097__A1 (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10097__B (.I(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10098__A1 (.I(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10098__A2 (.I(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10098__B1 (.I(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10098__B2 (.I(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__A2 (.I(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__B1 (.I(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10100__A1 (.I(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10100__A3 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10101__A1 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10101__B2 (.I(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10102__A1 (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10102__A2 (.I(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10103__A1 (.I(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10103__A2 (.I(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10105__B (.I(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10106__A1 (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10106__B (.I(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10107__A1 (.I(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10108__I0 (.I(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10108__S (.I(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10109__A1 (.I(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10109__A2 (.I(_04408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10109__B2 (.I(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10109__C (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__A1 (.I(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__B (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__B (.I(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10113__A1 (.I(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10113__A2 (.I(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10113__C (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10115__A2 (.I(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10115__B1 (.I(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10115__B2 (.I(\as2650.stack[11][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10116__A1 (.I(\as2650.stack[9][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10116__A2 (.I(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10116__B1 (.I(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__A1 (.I(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10118__A2 (.I(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10118__B1 (.I(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__A2 (.I(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__B1 (.I(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10120__A1 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10122__A2 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10122__B1 (.I(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10124__A2 (.I(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10124__B1 (.I(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10125__A1 (.I(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10126__I (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10127__I (.I(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10128__A2 (.I(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10128__B1 (.I(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10130__I (.I(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10131__A2 (.I(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10131__B1 (.I(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10132__A1 (.I(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10132__A2 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10133__A1 (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10133__B2 (.I(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__A2 (.I(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10135__A1 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10136__A1 (.I(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10138__A1 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10138__A2 (.I(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10140__A1 (.I(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10141__A1 (.I(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10141__A2 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10142__A1 (.I(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10142__A2 (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10143__A1 (.I(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10144__A1 (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10145__A1 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10146__B (.I(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10147__A2 (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10149__B2 (.I(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10151__A1 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10151__B (.I(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10153__A1 (.I(\as2650.instruction_args_latch[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10154__A2 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10155__A2 (.I(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10155__B1 (.I(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__A2 (.I(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__B1 (.I(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10157__A1 (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10158__A1 (.I(\as2650.stack[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10158__A2 (.I(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10158__B1 (.I(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10158__B2 (.I(\as2650.stack[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10159__A2 (.I(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10159__B1 (.I(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10160__A1 (.I(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10161__A1 (.I(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10162__A2 (.I(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10162__B1 (.I(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__A2 (.I(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__B1 (.I(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10164__A1 (.I(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10165__A1 (.I(\as2650.stack[13][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10165__A2 (.I(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10165__B1 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10166__A1 (.I(\as2650.stack[14][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10166__A2 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10166__B1 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10167__A1 (.I(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10168__A1 (.I(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10169__S (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10170__A2 (.I(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10171__A1 (.I(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__A1 (.I(\as2650.PC[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10173__B (.I(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10174__A1 (.I(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10174__A2 (.I(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10175__A1 (.I(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__A1 (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__B (.I(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10177__A1 (.I(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10177__B2 (.I(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__A1 (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__A2 (.I(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10180__A1 (.I(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10180__A2 (.I(_04408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10180__B2 (.I(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10182__A1 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10183__B (.I(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10185__B (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10187__A1 (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10187__A2 (.I(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10188__A1 (.I(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10188__A2 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10188__C (.I(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10190__A2 (.I(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10190__B1 (.I(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10191__I (.I(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10192__I (.I(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10193__B2 (.I(\as2650.stack[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10196__A1 (.I(\as2650.stack[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10196__A2 (.I(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10196__B1 (.I(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10197__A1 (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10197__A2 (.I(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10199__A2 (.I(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10199__B1 (.I(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10203__A2 (.I(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10203__B1 (.I(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10204__A1 (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10204__A2 (.I(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10205__A1 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10206__A1 (.I(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10207__A1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10207__A2 (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10208__A2 (.I(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10209__A1 (.I(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10210__A2 (.I(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10210__B2 (.I(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10211__I0 (.I(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10211__S (.I(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10212__I0 (.I(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__A1 (.I(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__A2 (.I(_04408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__B2 (.I(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10214__A1 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10215__B (.I(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10216__B (.I(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10218__A1 (.I(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10220__A1 (.I(\as2650.instruction_args_latch[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10220__A2 (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10220__B (.I(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10224__I (.I(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10225__I (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10227__I (.I(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10228__A1 (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10228__A2 (.I(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10229__A1 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10230__A2 (.I(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10231__A1 (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10232__I (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10234__A3 (.I(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10236__A1 (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10236__A2 (.I(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10237__A1 (.I(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10238__B (.I(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10239__A3 (.I(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10240__A1 (.I(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10241__I (.I(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10242__A1 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10242__A2 (.I(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10243__A1 (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10243__B (.I(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10243__C (.I(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10244__A4 (.I(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__I (.I(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10246__A1 (.I(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10247__A1 (.I(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10248__A1 (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10248__A2 (.I(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10250__A1 (.I(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10252__A1 (.I(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__B (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10260__A1 (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10260__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10263__A1 (.I(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10263__B (.I(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10264__A1 (.I(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10264__A2 (.I(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__A1 (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__A2 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10267__A1 (.I(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10267__A3 (.I(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10268__A1 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10271__A1 (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10272__A1 (.I(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10276__A1 (.I(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10276__A2 (.I(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10277__A1 (.I(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10278__A2 (.I(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10278__A3 (.I(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10282__I (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10284__A1 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10285__I (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__A1 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__B (.I(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10287__I (.I(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10289__I (.I(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__A1 (.I(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__A2 (.I(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__A1 (.I(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__A2 (.I(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10292__I (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10293__A1 (.I(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10294__A1 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10297__A1 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10297__A2 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10298__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10298__B (.I(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10300__A2 (.I(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10300__A3 (.I(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10302__I (.I(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10303__I (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10304__A1 (.I(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10307__A1 (.I(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10307__A2 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10308__A1 (.I(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10308__A2 (.I(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10313__A1 (.I(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10313__B1 (.I(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10313__B2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10315__A2 (.I(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10316__A1 (.I(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10317__A1 (.I(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10317__B2 (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10318__B (.I(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10320__A1 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10321__B (.I(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10324__S (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10325__A1 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__A1 (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__A1 (.I(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__A1 (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10329__A1 (.I(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__A1 (.I(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10331__B2 (.I(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__A1 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__A2 (.I(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10334__A1 (.I(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10334__A2 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10334__B (.I(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10336__A1 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10338__A1 (.I(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10338__A2 (.I(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10339__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10339__B (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__A1 (.I(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10341__A1 (.I(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10341__A2 (.I(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__A1 (.I(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__A2 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__A1 (.I(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__B1 (.I(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__B2 (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10344__A1 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10344__B2 (.I(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10345__B (.I(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10347__I (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10348__A1 (.I(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10348__A2 (.I(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10349__A1 (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10349__A2 (.I(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10350__I (.I(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10351__I (.I(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10352__A1 (.I(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10354__A1 (.I(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10354__A2 (.I(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10355__A1 (.I(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10355__A2 (.I(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10355__C (.I(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10356__A1 (.I(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10357__A1 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10359__A2 (.I(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10360__A1 (.I(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10360__A2 (.I(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10361__I (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10362__A1 (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10362__A2 (.I(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10362__B (.I(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10363__A1 (.I(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10364__A1 (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10366__A1 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10366__A2 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__A1 (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__A1 (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__A1 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__A2 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10372__A2 (.I(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10373__A1 (.I(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10379__A1 (.I(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10380__A1 (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10380__A2 (.I(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10380__A3 (.I(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10384__A1 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10386__A1 (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10387__A2 (.I(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10388__A1 (.I(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10388__A2 (.I(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10388__A3 (.I(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10390__A1 (.I(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10390__A2 (.I(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10391__A1 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10391__A2 (.I(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10391__A3 (.I(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10391__A4 (.I(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10392__A1 (.I(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10392__A2 (.I(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10392__A3 (.I(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10393__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10394__A1 (.I(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10396__A1 (.I(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10396__A2 (.I(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10396__A3 (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10399__A1 (.I(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10400__A1 (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10400__A2 (.I(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10400__A4 (.I(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10401__A1 (.I(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10402__A1 (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10402__A3 (.I(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10403__A3 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10404__A3 (.I(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10405__A1 (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__A1 (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__A2 (.I(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10407__A2 (.I(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10408__A1 (.I(\as2650.debug_psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10408__A3 (.I(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10410__I (.I(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10411__A1 (.I(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10413__A1 (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10413__A2 (.I(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10414__A1 (.I(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10414__A3 (.I(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10418__A1 (.I(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10418__A3 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10418__A4 (.I(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10420__A1 (.I(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10420__A2 (.I(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10420__A3 (.I(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10421__A1 (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10421__A2 (.I(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10422__B (.I(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10424__A1 (.I(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10425__A1 (.I(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10425__C (.I(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10426__A1 (.I(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10426__A2 (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10426__B1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10427__A1 (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10427__A2 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10428__A2 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10429__A1 (.I(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10429__A2 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__A1 (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10431__A1 (.I(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10431__A2 (.I(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10432__A2 (.I(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10433__A1 (.I(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10433__B1 (.I(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10433__B2 (.I(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__A1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__A2 (.I(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__B1 (.I(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__B2 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10435__A1 (.I(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10435__B1 (.I(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10436__A1 (.I(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10436__A2 (.I(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10437__A1 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10437__A2 (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10441__A1 (.I(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10441__A2 (.I(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10441__B1 (.I(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10441__B2 (.I(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10445__A1 (.I(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10445__A2 (.I(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10447__A1 (.I(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10448__B (.I(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10449__A3 (.I(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10450__A1 (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10453__A1 (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10453__A2 (.I(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10455__A1 (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10455__A2 (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10458__A1 (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10458__A2 (.I(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10459__A1 (.I(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10459__A2 (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10463__A1 (.I(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10464__A1 (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10465__A1 (.I(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10465__A2 (.I(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10465__B2 (.I(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10466__A1 (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10468__A1 (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10472__A2 (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10472__A3 (.I(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10472__A4 (.I(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10473__A1 (.I(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10473__A2 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10484__A1 (.I(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10485__A1 (.I(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10488__A1 (.I(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10489__A1 (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10492__A1 (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10492__A2 (.I(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10493__A1 (.I(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10493__A2 (.I(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10496__A2 (.I(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10498__A1 (.I(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10499__A1 (.I(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10500__A1 (.I(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10502__A1 (.I(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10505__A1 (.I(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10506__A1 (.I(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10511__A2 (.I(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10512__A1 (.I(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10513__A1 (.I(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10521__B (.I(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10527__A1 (.I(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10528__A2 (.I(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10531__A1 (.I(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10531__A2 (.I(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10533__A2 (.I(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10539__A1 (.I(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10539__A2 (.I(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10551__A1 (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10551__A2 (.I(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10552__A1 (.I(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10553__A1 (.I(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10557__A1 (.I(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10558__A1 (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10558__A3 (.I(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10558__A4 (.I(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10562__A1 (.I(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10579__A1 (.I(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10580__A2 (.I(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10587__A2 (.I(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10589__A2 (.I(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10592__A2 (.I(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10593__A1 (.I(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10597__A1 (.I(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10597__A2 (.I(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10609__A2 (.I(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10610__A2 (.I(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10616__A2 (.I(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10623__A3 (.I(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10624__B1 (.I(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10624__B2 (.I(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10626__A1 (.I(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10633__A1 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10634__A1 (.I(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10645__A2 (.I(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10646__A1 (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10655__A2 (.I(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10655__A3 (.I(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10655__A4 (.I(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10658__A2 (.I(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10664__A1 (.I(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10664__A2 (.I(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10675__A1 (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10676__A2 (.I(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10685__A1 (.I(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10686__A1 (.I(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10686__A2 (.I(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10687__A2 (.I(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10688__A2 (.I(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10689__A2 (.I(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10701__A2 (.I(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10704__A4 (.I(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10705__A1 (.I(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10705__A2 (.I(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10705__B1 (.I(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10707__A1 (.I(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10720__A1 (.I(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10735__A1 (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10751__A1 (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10751__A2 (.I(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10751__B1 (.I(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10751__B2 (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10752__A1 (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10752__A2 (.I(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10754__A1 (.I(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10754__A2 (.I(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10755__A1 (.I(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10755__A2 (.I(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10755__A3 (.I(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10756__A2 (.I(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10756__A3 (.I(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10759__A1 (.I(_05052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10759__A2 (.I(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10760__A1 (.I(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10762__A1 (.I(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10762__B (.I(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10764__A1 (.I(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10764__A2 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10764__A3 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10765__I (.I(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__A1 (.I(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10770__A1 (.I(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10770__A2 (.I(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10771__A1 (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10771__A2 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10771__B (.I(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10772__I (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10773__A1 (.I(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__A1 (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__A2 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__B (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10776__A1 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10776__B (.I(_03240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10778__A1 (.I(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10779__A1 (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10779__B (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10780__A1 (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10781__A1 (.I(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10781__A2 (.I(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10781__B (.I(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10783__A1 (.I(\as2650.debug_psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10785__A1 (.I(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10785__A2 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10785__B (.I(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10786__A1 (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10786__A2 (.I(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10788__A1 (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10788__A2 (.I(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10789__A1 (.I(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10789__A2 (.I(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10790__A2 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10793__A1 (.I(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10793__A2 (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10795__A1 (.I(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10795__A2 (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10796__A2 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10796__B1 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10796__B2 (.I(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10796__C1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10796__C2 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10797__A1 (.I(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10797__A2 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10797__B1 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10798__A1 (.I(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10798__A2 (.I(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10798__B1 (.I(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10798__B2 (.I(_03240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10799__A1 (.I(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10799__A2 (.I(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10804__A1 (.I(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10804__A2 (.I(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10804__B1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10804__B2 (.I(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10805__A2 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10805__B1 (.I(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10805__B2 (.I(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10806__A1 (.I(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10806__A2 (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10807__A2 (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10807__B1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10810__A1 (.I(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10810__A2 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10811__A2 (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10812__A1 (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10812__A2 (.I(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10813__A1 (.I(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10813__A2 (.I(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10814__I (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10815__A1 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10815__B1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10815__B2 (.I(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10816__A1 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10816__A2 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10817__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10817__A2 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10819__A1 (.I(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10819__A2 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10821__A2 (.I(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10822__A1 (.I(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10822__A2 (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10826__A1 (.I(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10826__A2 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10826__B1 (.I(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10826__B2 (.I(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10827__A1 (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10827__A2 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10829__A1 (.I(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10829__A2 (.I(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10829__A3 (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10830__A1 (.I(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10833__A1 (.I(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10833__A2 (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10834__A1 (.I(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10837__A1 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10838__A1 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10838__C (.I(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10840__C (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10841__A1 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10842__A2 (.I(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10843__A1 (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10845__A1 (.I(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10845__A2 (.I(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10846__A1 (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10846__A2 (.I(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10847__A1 (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10850__A2 (.I(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10851__A1 (.I(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10851__B1 (.I(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10851__B2 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10855__A1 (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10856__A2 (.I(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10856__B (.I(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10857__A1 (.I(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10857__A2 (.I(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10858__A2 (.I(_05052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10858__B2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10859__A1 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10861__A2 (.I(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10862__A1 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10864__A1 (.I(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10866__A1 (.I(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10867__A1 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10869__A1 (.I(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10870__A1 (.I(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10871__A1 (.I(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10871__A2 (.I(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10871__B (.I(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10872__A1 (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10872__B (.I(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10873__A1 (.I(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10874__A1 (.I(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10874__A2 (.I(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10875__A1 (.I(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10875__A2 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10876__A1 (.I(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10877__A1 (.I(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10878__A2 (.I(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10879__A1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10879__A2 (.I(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10880__A1 (.I(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10881__I (.I(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10883__I (.I(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10884__A1 (.I(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10885__A1 (.I(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10887__A1 (.I(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10888__A1 (.I(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10888__A2 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10888__B (.I(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10889__A1 (.I(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10889__A2 (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10891__A1 (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10892__A1 (.I(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10893__I (.I(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10895__A1 (.I(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10895__A2 (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10896__A1 (.I(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10896__A2 (.I(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10897__A1 (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10897__A2 (.I(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10898__A3 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10899__A3 (.I(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10899__B (.I(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10900__A1 (.I(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10901__A1 (.I(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10901__B (.I(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10902__I (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10903__A1 (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10904__A1 (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10905__A1 (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10906__B2 (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10907__I (.I(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10908__A1 (.I(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10910__A1 (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10910__A2 (.I(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10910__C (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10911__A1 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10911__A2 (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10914__A1 (.I(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10914__B (.I(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10916__A1 (.I(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10916__A2 (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10917__A1 (.I(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10917__A2 (.I(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__A1 (.I(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__A2 (.I(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10920__A1 (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10921__A1 (.I(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10922__A1 (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10923__A1 (.I(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10924__A1 (.I(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10926__B (.I(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10927__A1 (.I(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10928__A1 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10929__C (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10930__A1 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10930__B (.I(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10932__A1 (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10932__A2 (.I(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10933__A1 (.I(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10933__A2 (.I(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10935__A3 (.I(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10936__A1 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10936__A2 (.I(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10938__A1 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10940__A1 (.I(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10940__B (.I(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10943__A1 (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10943__A2 (.I(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10944__A1 (.I(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10944__A2 (.I(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10945__A1 (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10946__A2 (.I(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10946__B (.I(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10948__I (.I(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10950__B (.I(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__A1 (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__B2 (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10953__A1 (.I(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10954__I (.I(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10955__A1 (.I(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10955__A2 (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10955__B (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10956__A1 (.I(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10957__B2 (.I(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10957__C (.I(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10958__I (.I(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10959__A1 (.I(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10959__A2 (.I(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10959__B2 (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10960__B2 (.I(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10961__A1 (.I(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10961__A2 (.I(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10961__A3 (.I(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10962__A1 (.I(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10962__B1 (.I(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10963__A1 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10963__A2 (.I(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10964__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10964__B (.I(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10965__A2 (.I(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10966__A1 (.I(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10967__A1 (.I(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10967__A2 (.I(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10967__C (.I(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10968__A1 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10968__B2 (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10970__A1 (.I(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10971__A1 (.I(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10971__A2 (.I(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10972__A1 (.I(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10972__A2 (.I(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10972__B (.I(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10973__C (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10974__A1 (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10974__B2 (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10976__A1 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10977__A1 (.I(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10977__A2 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10977__C (.I(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10978__I (.I(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10979__C (.I(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10980__A1 (.I(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10981__I (.I(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10988__I (.I(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10989__I0 (.I(\as2650.trap ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10998__A1 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10998__A3 (.I(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10999__B2 (.I(\as2650.trap ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11000__A1 (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11001__I (.I(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11004__B (.I(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11005__A1 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11006__B (.I(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11007__A1 (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11011__A1 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11013__A1 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__A1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__A1 (.I(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11019__B (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11020__A1 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11021__B (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11022__A1 (.I(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11023__A1 (.I(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11023__A2 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11023__B (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11025__I (.I(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11027__A2 (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11028__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11028__C (.I(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11029__A2 (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11030__A1 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11030__C (.I(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11031__A1 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11031__A2 (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11032__A1 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11032__C (.I(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11035__I (.I(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11036__A1 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11039__A1 (.I(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11040__A1 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11041__A1 (.I(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11042__A1 (.I(\as2650.ext_io_addr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11043__A1 (.I(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11044__A1 (.I(\as2650.ext_io_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11045__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11045__C (.I(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11046__A1 (.I(\as2650.io_bus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11047__A1 (.I(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11050__A2 (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11051__A3 (.I(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11051__A4 (.I(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11052__A1 (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11052__A2 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11052__A3 (.I(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11053__A1 (.I(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11053__A2 (.I(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11053__B2 (.I(_05331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11054__A2 (.I(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11055__A1 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11056__A1 (.I(_05333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11057__I (.I(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11058__A1 (.I(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11059__A1 (.I(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11059__A2 (.I(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11060__I (.I(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11062__A1 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11064__I (.I(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11065__I (.I(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11066__A1 (.I(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11066__A2 (.I(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11066__B (.I(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11066__C (.I(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11067__I (.I(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11068__A1 (.I(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11069__A1 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11070__I (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11071__A1 (.I(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11071__B2 (.I(\as2650.regs[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11072__A1 (.I(_03035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11073__I (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11074__A1 (.I(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11075__A1 (.I(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11076__I (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11077__A1 (.I(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11078__A1 (.I(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11079__I (.I(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11080__I (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11081__I (.I(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11082__I (.I(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__A1 (.I(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11084__A1 (.I(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11085__I (.I(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11086__A1 (.I(_05358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11087__A1 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11088__I (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11089__A1 (.I(_05360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11089__B2 (.I(\as2650.regs[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11091__I (.I(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11092__A1 (.I(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11092__B2 (.I(\as2650.regs[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11094__A2 (.I(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11094__A3 (.I(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11096__A2 (.I(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11097__I (.I(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__A1 (.I(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11099__A1 (.I(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11099__A2 (.I(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11101__A1 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11102__A1 (.I(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11104__A1 (.I(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11104__A2 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11105__A2 (.I(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11105__A3 (.I(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11107__A2 (.I(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11113__A1 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11114__A2 (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11115__A1 (.I(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11116__A1 (.I(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11116__A2 (.I(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11116__A3 (.I(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11119__A1 (.I(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11119__A2 (.I(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11120__A2 (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11126__A2 (.I(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11127__I (.I(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11130__A1 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11136__I (.I(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11137__I (.I(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11138__A1 (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11139__A1 (.I(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11142__A1 (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11142__A2 (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11145__A1 (.I(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11147__A1 (.I(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11150__A1 (.I(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11155__I (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11157__A3 (.I(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11158__A1 (.I(_05427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11158__A2 (.I(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11160__A1 (.I(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11160__B1 (.I(_05429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11160__B2 (.I(\as2650.regs[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11162__A1 (.I(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11163__I (.I(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11164__A1 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11164__A2 (.I(_05427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11164__C (.I(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11170__A1 (.I(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11171__A1 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11171__A2 (.I(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11171__A3 (.I(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11174__A1 (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11178__A1 (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11180__A1 (.I(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11181__A1 (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11183__A2 (.I(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11186__A1 (.I(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11186__A2 (.I(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11186__B1 (.I(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11190__A1 (.I(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11193__A1 (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11193__A2 (.I(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11194__A1 (.I(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11198__A1 (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11199__A1 (.I(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11202__A1 (.I(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11203__A2 (.I(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11204__A1 (.I(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__A1 (.I(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__B1 (.I(_05429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__B2 (.I(\as2650.regs[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11209__A1 (.I(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11210__A1 (.I(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11211__A1 (.I(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11215__A1 (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11216__A1 (.I(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11218__A1 (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11219__A2 (.I(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11220__A1 (.I(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11221__A1 (.I(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11221__B1 (.I(_05429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11221__B2 (.I(\as2650.regs[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11224__A1 (.I(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11226__I (.I(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11227__A1 (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11228__A1 (.I(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11231__A1 (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11232__A1 (.I(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11233__A1 (.I(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11234__A1 (.I(\as2650.regs[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11235__A1 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11236__A2 (.I(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11237__A1 (.I(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11237__B1 (.I(_05429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11240__A1 (.I(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11242__A1 (.I(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11243__A1 (.I(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11245__A1 (.I(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11246__A1 (.I(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11247__A1 (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11248__A1 (.I(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11250__A1 (.I(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11251__A1 (.I(_05358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11251__A2 (.I(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11251__B1 (.I(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11253__A1 (.I(\as2650.regs[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11254__A1 (.I(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11255__A1 (.I(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11256__A1 (.I(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11258__A1 (.I(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11259__A1 (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11261__A1 (.I(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11262__A1 (.I(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11263__A1 (.I(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11265__A1 (.I(_05360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11265__A2 (.I(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11265__B1 (.I(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11265__B2 (.I(\as2650.regs[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11267__A1 (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11268__A1 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11269__A1 (.I(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11270__A1 (.I(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11271__A1 (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11273__A1 (.I(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11274__A1 (.I(\as2650.regs[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11275__A1 (.I(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11275__B2 (.I(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11276__A1 (.I(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11277__A1 (.I(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11277__A2 (.I(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11277__B1 (.I(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11277__B2 (.I(\as2650.regs[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11279__A2 (.I(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11280__A1 (.I(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11280__A2 (.I(_05541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11281__I (.I(_05542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11282__I (.I(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11284__I (.I(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11289__A1 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11291__A1 (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11292__A1 (.I(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11294__I (.I(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11295__I (.I(_05542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11296__A1 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11296__A3 (.I(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11296__A4 (.I(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11298__A1 (.I(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11298__B1 (.I(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11298__C2 (.I(\as2650.regs[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11299__A1 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11301__A1 (.I(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11303__A1 (.I(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11304__A1 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11306__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11306__B1 (.I(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11306__C2 (.I(\as2650.regs[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11307__A1 (.I(_03035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11308__I (.I(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11311__A1 (.I(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11313__A1 (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11314__A1 (.I(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11315__A1 (.I(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11317__A1 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11317__B2 (.I(\as2650.regs[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11317__C (.I(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11318__A1 (.I(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11320__A1 (.I(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11321__A1 (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11323__A1 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11323__B1 (.I(_05581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11324__A1 (.I(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11325__I (.I(_05542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11326__A1 (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11327__A1 (.I(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11331__A1 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11331__C (.I(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11332__A1 (.I(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11333__A1 (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11334__A1 (.I(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11338__A1 (.I(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11338__C (.I(_05594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11339__A1 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11340__A1 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11341__A1 (.I(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11345__A1 (.I(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11345__B2 (.I(\as2650.regs[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11345__C (.I(_05600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11347__A1 (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11348__A1 (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11349__A1 (.I(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11349__A2 (.I(_05052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11350__A1 (.I(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11350__B1 (.I(_05604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11350__C2 (.I(\as2650.regs[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11352__A1 (.I(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11352__A2 (.I(_05541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11353__I (.I(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11355__I (.I(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11356__A1 (.I(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11356__A2 (.I(_05541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11356__B (.I(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11356__C (.I(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11357__I (.I(_05610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11358__A1 (.I(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__A1 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11360__A1 (.I(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11361__A1 (.I(_03035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11362__A1 (.I(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11363__A1 (.I(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11364__A1 (.I(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11365__A1 (.I(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11366__I (.I(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11367__I (.I(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11368__I (.I(_05610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11369__A1 (.I(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11369__B2 (.I(\as2650.regs[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11370__A1 (.I(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11371__A1 (.I(_05358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11371__B2 (.I(\as2650.regs[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11372__A1 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11373__A1 (.I(_05360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11373__B2 (.I(\as2650.regs[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11375__A1 (.I(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11375__B2 (.I(\as2650.regs[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11377__A3 (.I(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11378__I (.I(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11383__I (.I(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11384__A1 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11386__A1 (.I(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11386__B2 (.I(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11386__C1 (.I(\as2650.regs[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11387__A1 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11388__A1 (.I(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11388__B2 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11388__C1 (.I(\as2650.regs[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11389__A1 (.I(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11392__A1 (.I(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11394__A1 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11394__B2 (.I(\as2650.regs[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11395__A1 (.I(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11396__A1 (.I(_05581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11396__B2 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11396__C1 (.I(\as2650.regs[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11397__A1 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11398__I (.I(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11400__A1 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11400__B2 (.I(\as2650.regs[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11401__A1 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11403__A1 (.I(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11404__A1 (.I(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11406__A1 (.I(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11406__B2 (.I(\as2650.regs[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11407__A1 (.I(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11408__A1 (.I(_05604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11408__B2 (.I(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11408__C1 (.I(\as2650.regs[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11409__A1 (.I(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11410__A3 (.I(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11411__I (.I(_05648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11413__I (.I(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11414__I (.I(_05648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11415__A1 (.I(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11415__A2 (.I(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11417__A1 (.I(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11418__A1 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11419__A1 (.I(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11419__B2 (.I(\as2650.regs[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11420__A1 (.I(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11421__A1 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11422__A1 (.I(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11423__A1 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11423__B2 (.I(\as2650.regs[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11424__A1 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11425__I (.I(_05648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11426__I (.I(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11428__A1 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11428__B2 (.I(\as2650.regs[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11429__A1 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11430__A1 (.I(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11430__B2 (.I(\as2650.regs[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11431__A1 (.I(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11432__A1 (.I(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11432__B2 (.I(\as2650.regs[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11433__A1 (.I(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11434__A1 (.I(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11434__B2 (.I(\as2650.regs[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11435__A1 (.I(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11437__A1 (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11437__A2 (.I(_05541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11441__A2 (.I(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11441__B2 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11442__A1 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11442__A2 (.I(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11442__A3 (.I(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11442__A4 (.I(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11444__A1 (.I(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11444__A2 (.I(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11447__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11448__I (.I(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11449__A1 (.I(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11451__A1 (.I(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11451__B1 (.I(_05680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11451__B2 (.I(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11453__A1 (.I(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11453__A2 (.I(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11455__A2 (.I(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11456__A1 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11456__A2 (.I(_05682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11456__B2 (.I(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11458__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11458__A2 (.I(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11463__A1 (.I(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11463__A2 (.I(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11464__A1 (.I(\as2650.regs[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11465__A1 (.I(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11465__B2 (.I(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11467__A1 (.I(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11467__B1 (.I(_05680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11469__A1 (.I(\as2650.regs[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11470__A1 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11470__B2 (.I(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11472__A1 (.I(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11472__B1 (.I(_05680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11474__A1 (.I(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11474__A2 (.I(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11474__B2 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11475__A1 (.I(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11476__I (.I(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11477__A1 (.I(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11477__B1 (.I(_05680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11477__B2 (.I(\as2650.regs[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11479__A1 (.I(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11479__A2 (.I(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11479__B2 (.I(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11482__A1 (.I(_05358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11484__A1 (.I(\as2650.regs[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11485__A1 (.I(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11488__A1 (.I(_05360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11488__B2 (.I(\as2650.regs[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11490__A1 (.I(\as2650.regs[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11491__A1 (.I(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11491__B2 (.I(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11493__A1 (.I(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11493__B2 (.I(\as2650.regs[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11495__A1 (.I(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11496__I (.I(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11497__S (.I(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11499__S (.I(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11501__S (.I(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11503__S (.I(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11505__I (.I(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11506__S (.I(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11508__I1 (.I(\as2650.stack[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11508__S (.I(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11510__I1 (.I(\as2650.stack[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11510__S (.I(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11512__S (.I(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11514__I (.I(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11515__I0 (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11517__I0 (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11519__I0 (.I(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11519__I1 (.I(\as2650.stack[9][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11521__I0 (.I(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11523__I (.I(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11524__S (.I(_05733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11526__S (.I(_05733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11528__S (.I(_05733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11530__S (.I(_05733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11532__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11568__CLK (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11771__CLK (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11842__CLK (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11874__D (.I(_00342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11876__D (.I(_00344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11908__CLK (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11909__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11913__CLK (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11931__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11932__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11933__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11934__CLK (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11935__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11982__CLK (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11985__CLK (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11987__D (.I(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11990__D (.I(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11991__D (.I(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11993__CLK (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11993__D (.I(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11994__D (.I(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11996__D (.I(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11998__CLK (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11998__D (.I(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11999__D (.I(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12000__CLK (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12004__D (.I(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12005__CLK (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12045__CLK (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12097__CLK (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12110__CLK (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12157__I (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12158__I (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12159__I (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12160__I (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12161__I (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12162__I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12163__I (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12164__I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_0__f_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_10__f_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_11__f_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_12__f_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_13__f_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_14__f_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_15__f_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_1__f_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_2__f_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_3__f_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_4__f_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_5__f_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_6__f_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_7__f_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_8__f_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_9__f_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_101_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_102_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_103_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_104_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_105_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_106_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_107_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_108_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_109_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_110_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_111_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_112_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_113_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_114_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_115_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_116_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_117_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_118_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_119_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_120_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_121_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_122_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_123_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_124_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_125_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_126_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_127_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_128_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_130_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_131_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_132_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_133_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_134_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_135_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_136_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_137_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_138_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_139_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_140_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_141_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_142_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_143_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_144_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_145_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_146_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_147_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_148_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_149_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_150_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_152_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_153_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_154_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_155_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_156_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_157_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_158_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_159_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_160_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_161_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_162_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_163_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_164_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_165_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_166_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_167_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_64_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_70_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_72_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_73_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_75_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_78_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_79_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_80_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_81_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_82_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_83_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_85_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_87_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_88_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_89_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_90_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_91_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_92_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_93_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_94_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_95_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_96_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_97_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_98_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_99_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout250_I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout251_I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold100_I (.I(wbs_dat_i[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold101_I (.I(wbs_dat_i[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold102_I (.I(wbs_dat_i[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold103_I (.I(wbs_dat_i[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold104_I (.I(wbs_dat_i[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold105_I (.I(wbs_dat_i[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold106_I (.I(wbs_dat_i[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold107_I (.I(wbs_dat_i[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold108_I (.I(wbs_dat_i[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold109_I (.I(wbs_dat_i[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold110_I (.I(wbs_dat_i[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold111_I (.I(wbs_dat_i[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold112_I (.I(wbs_dat_i[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold113_I (.I(wbs_dat_i[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold114_I (.I(wbs_dat_i[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold115_I (.I(wbs_dat_i[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold116_I (.I(wbs_dat_i[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold117_I (.I(wbs_dat_i[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold118_I (.I(wbs_dat_i[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold119_I (.I(wbs_dat_i[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold120_I (.I(wbs_adr_i[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold12_I (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold20_I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold30_I (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold38_I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold42_I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold50_I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold53_I (.I(wbs_adr_i[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold54_I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold64_I (.I(wbs_adr_i[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold67_I (.I(wbs_dat_i[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold85_I (.I(wbs_cyc_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold86_I (.I(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold87_I (.I(wbs_dat_i[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold88_I (.I(wbs_dat_i[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold89_I (.I(wbs_dat_i[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold90_I (.I(wbs_dat_i[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold91_I (.I(wbs_dat_i[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold92_I (.I(wbs_dat_i[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold93_I (.I(wbs_dat_i[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold94_I (.I(wbs_dat_i[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold95_I (.I(wbs_dat_i[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold96_I (.I(wbs_dat_i[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold97_I (.I(wbs_adr_i[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold98_I (.I(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold99_I (.I(wbs_dat_i[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(bus_in_serial_ports[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(bus_in_serial_ports[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(bus_in_serial_ports[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(bus_in_serial_ports[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(bus_in_serial_ports[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(bus_in_serial_ports[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(bus_in_serial_ports[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(bus_in_timers[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(bus_in_timers[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(bus_in_timers[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(bus_in_gpios[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(bus_in_timers[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(bus_in_timers[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(bus_in_timers[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(bus_in_timers[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(bus_in_timers[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(bus_in_gpios[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(irqs[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(irqs[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(irqs[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(irqs[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(irqs[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(bus_in_gpios[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(irqs[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(irqs[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(rom_bus_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(rom_bus_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(rom_bus_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(rom_bus_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(rom_bus_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(rom_bus_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(rom_bus_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(rom_bus_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(bus_in_gpios[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(wb_rst_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(bus_in_gpios[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(bus_in_gpios[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(bus_in_gpios[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input88_I (.I(wbs_stb_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input89_I (.I(wbs_we_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(bus_in_gpios[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(bus_in_serial_ports[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap252_I (.I(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output100_I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output101_I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output102_I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output103_I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output104_I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output105_I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output106_I (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output107_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output108_I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output109_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output110_I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output111_I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output112_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output113_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output114_I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output115_I (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output116_I (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output117_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output118_I (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output119_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output120_I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output121_I (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output123_I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output126_I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output129_I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output130_I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output142_I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output143_I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output144_I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output148_I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output154_I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output155_I (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output156_I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output157_I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output158_I (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output159_I (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output160_I (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output161_I (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output162_I (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output163_I (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output164_I (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output165_I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output166_I (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output167_I (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output168_I (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output169_I (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output170_I (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output171_I (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output172_I (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output173_I (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output174_I (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output175_I (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output176_I (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output177_I (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output178_I (.I(net178));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output179_I (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output180_I (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output181_I (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output182_I (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output183_I (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output184_I (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output187_I (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output188_I (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output189_I (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output190_I (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output191_I (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output192_I (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output193_I (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output194_I (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output195_I (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output196_I (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output197_I (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output198_I (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output199_I (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output200_I (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output201_I (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output202_I (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output203_I (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output204_I (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output205_I (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output206_I (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output236_I (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output237_I (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output239_I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output240_I (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output90_I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output91_I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output92_I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output93_I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output94_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output95_I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output96_I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output97_I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output98_I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output99_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer1_I (.I(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer3_I (.I(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer8_I (.I(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_157_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_157_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_163_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_163_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_165_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_165_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_167_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_168_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_168_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_168_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_998 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Left_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Left_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Left_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Left_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Left_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Left_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Left_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Left_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Left_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Left_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Left_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Left_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Left_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Left_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Left_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Left_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Left_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Left_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Left_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Left_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Left_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Left_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Left_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Left_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Left_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Left_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Left_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Left_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Left_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Left_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Left_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Left_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Left_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Left_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Left_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Left_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Left_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Left_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Left_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Left_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Left_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Left_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Left_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Left_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Left_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_Left_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_Right_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_Left_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_Right_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_Left_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_Right_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_Left_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_Right_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_Left_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_Right_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_Left_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_Right_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_Left_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_Right_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_Left_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_Right_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_Left_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_Right_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_Left_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_Right_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_Left_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_Right_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_Left_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_Right_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_Left_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_Right_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_Left_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_Right_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_Left_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_Right_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_Left_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_Right_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_Left_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_Right_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_Left_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_Right_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_Left_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_Right_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_Left_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_Right_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_Left_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_Right_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_Left_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_Right_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_Left_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_Right_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_Left_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_Right_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_Left_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_Right_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Left_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Left_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Left_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Left_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Left_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Left_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Left_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Left_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Left_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Left_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Left_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Left_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Left_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Left_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Left_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Left_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Left_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Left_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Left_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Left_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Left_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Left_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Left_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Left_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Left_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Left_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Left_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Left_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Left_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_615 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05738_ (.I(\as2650.debug_psl[4] ),
    .Z(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05739_ (.I(_00579_),
    .Z(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05740_ (.I(_00580_),
    .Z(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05741_ (.I(_00581_),
    .Z(_00582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05742_ (.I(_00582_),
    .Z(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05743_ (.I0(\as2650.regs[1][7] ),
    .I1(\as2650.regs[5][7] ),
    .S(_00583_),
    .Z(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05744_ (.I(_00584_),
    .Z(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05745_ (.I(_00585_),
    .Z(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05746_ (.I(_00586_),
    .Z(_00587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05747_ (.I(_00587_),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05748_ (.I0(\as2650.regs[1][6] ),
    .I1(\as2650.regs[5][6] ),
    .S(_00583_),
    .Z(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05749_ (.I(_00588_),
    .Z(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _05750_ (.I(_00589_),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05751_ (.I(_00579_),
    .Z(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05752_ (.I0(\as2650.regs[1][5] ),
    .I1(\as2650.regs[5][5] ),
    .S(_00590_),
    .Z(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05753_ (.I(_00591_),
    .Z(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05754_ (.I(_00592_),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05755_ (.I(_00579_),
    .Z(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05756_ (.I0(\as2650.regs[1][4] ),
    .I1(\as2650.regs[5][4] ),
    .S(_00593_),
    .Z(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05757_ (.I(_00594_),
    .Z(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05758_ (.I(_00595_),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05759_ (.I0(\as2650.regs[1][3] ),
    .I1(\as2650.regs[5][3] ),
    .S(_00581_),
    .Z(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05760_ (.I(_00596_),
    .Z(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05761_ (.I(_00597_),
    .Z(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05762_ (.I(_00598_),
    .Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05763_ (.I0(\as2650.regs[1][2] ),
    .I1(\as2650.regs[5][2] ),
    .S(_00582_),
    .Z(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05764_ (.I(_00599_),
    .Z(_00600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05765_ (.I(_00600_),
    .Z(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05766_ (.I(_00601_),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05767_ (.I0(\as2650.regs[1][1] ),
    .I1(\as2650.regs[5][1] ),
    .S(_00581_),
    .Z(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05768_ (.I(_00602_),
    .Z(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05769_ (.I(_00603_),
    .Z(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05770_ (.I(_00604_),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05771_ (.I0(\as2650.regs[1][0] ),
    .I1(\as2650.regs[5][0] ),
    .S(_00582_),
    .Z(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05772_ (.I(_00605_),
    .Z(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05773_ (.I(_00606_),
    .Z(_00607_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05774_ (.I(_00607_),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05775_ (.A1(_00583_),
    .A2(\as2650.regs[4][7] ),
    .ZN(_00608_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05776_ (.I(\as2650.debug_psl[4] ),
    .ZN(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05777_ (.I(_00609_),
    .Z(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05778_ (.I(_00610_),
    .Z(_00611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05779_ (.I(_00611_),
    .Z(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05780_ (.A1(_00612_),
    .A2(\as2650.regs[0][7] ),
    .ZN(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05781_ (.A1(_00608_),
    .A2(_00613_),
    .Z(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05782_ (.I(_00614_),
    .ZN(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05783_ (.I(_00615_),
    .Z(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05784_ (.I(_00616_),
    .Z(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05785_ (.I(_00617_),
    .Z(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05786_ (.I(_00618_),
    .Z(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05787_ (.I(_00619_),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05788_ (.I0(\as2650.regs[0][6] ),
    .I1(\as2650.regs[4][6] ),
    .S(_00582_),
    .Z(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05789_ (.I(_00620_),
    .Z(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05790_ (.I(_00621_),
    .Z(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _05791_ (.I(_00622_),
    .Z(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05792_ (.I(_00623_),
    .Z(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05793_ (.I(_00624_),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05794_ (.A1(_00611_),
    .A2(\as2650.regs[0][5] ),
    .ZN(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05795_ (.A1(_00590_),
    .A2(\as2650.regs[4][5] ),
    .ZN(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _05796_ (.A1(_00625_),
    .A2(_00626_),
    .Z(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05797_ (.I(_00627_),
    .ZN(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05798_ (.I(_00628_),
    .Z(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05799_ (.I(_00629_),
    .Z(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05800_ (.I(_00630_),
    .Z(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05801_ (.I(_00631_),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05802_ (.I(\as2650.regs[4][4] ),
    .ZN(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05803_ (.A1(_00580_),
    .A2(_00632_),
    .ZN(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05804_ (.A1(_00590_),
    .A2(\as2650.regs[0][4] ),
    .B(_00633_),
    .ZN(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05805_ (.I(_00634_),
    .ZN(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05806_ (.I(_00635_),
    .Z(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05807_ (.I(_00636_),
    .Z(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05808_ (.I(_00637_),
    .Z(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05809_ (.I(_00638_),
    .Z(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05810_ (.I(_00639_),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05811_ (.I(\as2650.cycle[3] ),
    .Z(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05812_ (.I(_00640_),
    .ZN(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05813_ (.I(\as2650.cycle[1] ),
    .Z(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05814_ (.I(_00642_),
    .Z(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05815_ (.I(_00643_),
    .ZN(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05816_ (.I(_00644_),
    .Z(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05817_ (.I(\as2650.cycle[2] ),
    .Z(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05818_ (.A1(_00645_),
    .A2(_00646_),
    .ZN(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05819_ (.A1(_00641_),
    .A2(_00647_),
    .ZN(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05820_ (.I(_00648_),
    .Z(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05821_ (.I(_00649_),
    .Z(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05822_ (.I(_00650_),
    .Z(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _05823_ (.I(\as2650.relative_cyc ),
    .ZN(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05824_ (.I(\as2650.cycle[0] ),
    .Z(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05825_ (.I(_00653_),
    .Z(_00654_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05826_ (.A1(_00646_),
    .A2(_00640_),
    .ZN(_00655_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _05827_ (.A1(_00654_),
    .A2(_00643_),
    .A3(_00655_),
    .ZN(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05828_ (.I(_00656_),
    .Z(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05829_ (.I(\as2650.indirect_cyc ),
    .Z(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05830_ (.A1(_00658_),
    .A2(_00648_),
    .ZN(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _05831_ (.A1(_00652_),
    .A2(_00657_),
    .A3(_00659_),
    .ZN(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05832_ (.A1(\as2650.indexed_cyc[1] ),
    .A2(\as2650.indexed_cyc[0] ),
    .ZN(_00661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05833_ (.A1(\as2650.wb_hidden_rom_enable ),
    .A2(\as2650.cpu_hidden_rom_enable ),
    .ZN(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05834_ (.I(_00662_),
    .Z(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05835_ (.I(_00663_),
    .Z(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05836_ (.I(\as2650.wb_hidden_rom_enable ),
    .Z(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05837_ (.I(_00665_),
    .Z(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05838_ (.I(_00666_),
    .Z(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05839_ (.I(\as2650.cpu_hidden_rom_enable ),
    .Z(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05840_ (.I(_00668_),
    .Z(_00669_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05841_ (.A1(_00667_),
    .A2(_00669_),
    .A3(net49),
    .Z(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _05842_ (.A1(\as2650.cycle[0] ),
    .A2(\as2650.cycle[1] ),
    .A3(\as2650.cycle[2] ),
    .A4(\as2650.cycle[3] ),
    .Z(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _05843_ (.I(_00671_),
    .Z(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05844_ (.I(_00672_),
    .Z(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05845_ (.I(_00673_),
    .Z(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05846_ (.A1(net28),
    .A2(_00664_),
    .B(_00670_),
    .C(_00674_),
    .ZN(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05847_ (.A1(_00653_),
    .A2(_00642_),
    .A3(\as2650.cycle[2] ),
    .A4(net302),
    .ZN(_00676_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05848_ (.I(net379),
    .Z(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05849_ (.A1(\as2650.insin[7] ),
    .A2(_00677_),
    .ZN(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05850_ (.A1(\as2650.insin[6] ),
    .A2(_00674_),
    .Z(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05851_ (.I(net48),
    .ZN(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05852_ (.I(_00662_),
    .ZN(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05853_ (.I(_00681_),
    .Z(_00682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05854_ (.I(_00682_),
    .Z(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _05855_ (.I(_00666_),
    .Z(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05856_ (.A1(_00684_),
    .A2(_00669_),
    .B(net27),
    .ZN(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05857_ (.A1(_00680_),
    .A2(_00683_),
    .B(_00685_),
    .C(_00674_),
    .ZN(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05858_ (.A1(_00675_),
    .A2(_00678_),
    .A3(_00679_),
    .A4(_00686_),
    .ZN(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05859_ (.I(_00673_),
    .Z(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05860_ (.A1(\as2650.insin[4] ),
    .A2(_00688_),
    .Z(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05861_ (.I(net46),
    .ZN(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05862_ (.I(_00668_),
    .Z(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05863_ (.A1(_00667_),
    .A2(_00691_),
    .B(net34),
    .ZN(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05864_ (.A1(_00690_),
    .A2(_00683_),
    .B(_00692_),
    .C(_00688_),
    .ZN(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05865_ (.A1(\as2650.insin[5] ),
    .A2(_00688_),
    .Z(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05866_ (.I(net47),
    .ZN(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05867_ (.A1(_00667_),
    .A2(_00691_),
    .B(net26),
    .ZN(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05868_ (.A1(_00695_),
    .A2(_00682_),
    .B(_00696_),
    .C(_00673_),
    .ZN(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _05869_ (.A1(_00689_),
    .A2(_00693_),
    .A3(_00694_),
    .A4(_00697_),
    .Z(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05870_ (.I(_00673_),
    .Z(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05871_ (.A1(\as2650.insin[7] ),
    .A2(_00699_),
    .Z(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05872_ (.I(net49),
    .ZN(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05873_ (.A1(_00684_),
    .A2(_00669_),
    .B(net28),
    .ZN(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05874_ (.A1(_00701_),
    .A2(_00683_),
    .B(_00702_),
    .C(_00688_),
    .ZN(_00703_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _05875_ (.A1(_00666_),
    .A2(_00668_),
    .A3(net48),
    .Z(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05876_ (.A1(net27),
    .A2(_00663_),
    .B(_00704_),
    .C(_00699_),
    .ZN(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05877_ (.A1(\as2650.insin[6] ),
    .A2(net379),
    .ZN(_00706_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05878_ (.A1(_00700_),
    .A2(_00703_),
    .A3(_00705_),
    .A4(_00706_),
    .ZN(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05879_ (.I(\as2650.extend ),
    .Z(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _05880_ (.A1(_00687_),
    .A2(_00698_),
    .A3(_00707_),
    .B(_00708_),
    .ZN(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _05881_ (.A1(_00666_),
    .A2(_00691_),
    .A3(net45),
    .Z(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05882_ (.A1(net33),
    .A2(_00663_),
    .B(_00710_),
    .C(_00699_),
    .ZN(_00711_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05883_ (.A1(\as2650.insin[3] ),
    .A2(net380),
    .ZN(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _05884_ (.A1(_00711_),
    .A2(_00712_),
    .Z(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05885_ (.I(_00699_),
    .Z(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05886_ (.I0(net32),
    .I1(net44),
    .S(_00682_),
    .Z(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05887_ (.A1(\as2650.insin[2] ),
    .A2(_00677_),
    .Z(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05888_ (.A1(_00714_),
    .A2(_00715_),
    .B(_00716_),
    .ZN(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _05889_ (.A1(\as2650.indirect_cyc ),
    .A2(_00713_),
    .A3(_00717_),
    .ZN(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _05890_ (.A1(_00667_),
    .A2(_00691_),
    .A3(net46),
    .Z(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05891_ (.A1(net34),
    .A2(_00663_),
    .B(_00719_),
    .C(_00674_),
    .ZN(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05892_ (.A1(\as2650.insin[4] ),
    .A2(_00677_),
    .ZN(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05893_ (.A1(_00720_),
    .A2(_00721_),
    .A3(_00711_),
    .A4(_00712_),
    .ZN(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05894_ (.I(\as2650.instruction_args_latch[13] ),
    .Z(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05895_ (.A1(_00723_),
    .A2(\as2650.instruction_args_latch[14] ),
    .ZN(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05896_ (.I(\as2650.extend ),
    .ZN(_00725_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05897_ (.A1(_00722_),
    .A2(_00724_),
    .B(_00725_),
    .ZN(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _05898_ (.A1(_00709_),
    .A2(_00718_),
    .A3(_00726_),
    .ZN(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05899_ (.A1(_00656_),
    .A2(_00661_),
    .B(_00727_),
    .ZN(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05900_ (.A1(_00660_),
    .A2(_00728_),
    .Z(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05901_ (.I(_00729_),
    .Z(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _05902_ (.I(\as2650.instruction_args_latch[14] ),
    .ZN(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05903_ (.I(\as2650.indexed_cyc[1] ),
    .ZN(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05904_ (.A1(\as2650.indexed_cyc[0] ),
    .A2(_00731_),
    .B(_00732_),
    .ZN(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05905_ (.A1(_00708_),
    .A2(_00733_),
    .ZN(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05906_ (.I(\as2650.instruction_args_latch[13] ),
    .ZN(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05907_ (.I(\as2650.indexed_cyc[0] ),
    .ZN(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05908_ (.A1(\as2650.indexed_cyc[1] ),
    .A2(_00735_),
    .B(_00736_),
    .ZN(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _05909_ (.A1(_00734_),
    .A2(_00737_),
    .ZN(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05910_ (.I(_00738_),
    .Z(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _05911_ (.A1(_00665_),
    .A2(net42),
    .A3(\as2650.cpu_hidden_rom_enable ),
    .Z(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05912_ (.A1(net30),
    .A2(_00662_),
    .B(_00740_),
    .C(_00672_),
    .ZN(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05913_ (.I(_00741_),
    .Z(_00742_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05914_ (.A1(\as2650.insin[0] ),
    .A2(_00676_),
    .ZN(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05915_ (.I(_00743_),
    .Z(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05916_ (.A1(_00742_),
    .A2(_00744_),
    .ZN(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05917_ (.I(_00745_),
    .Z(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _05918_ (.A1(\as2650.insin[0] ),
    .A2(net297),
    .Z(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05919_ (.I(_00747_),
    .Z(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05920_ (.I(_00748_),
    .Z(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05921_ (.I(net42),
    .ZN(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05922_ (.A1(_00665_),
    .A2(\as2650.cpu_hidden_rom_enable ),
    .B(net30),
    .ZN(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05923_ (.A1(_00750_),
    .A2(_00681_),
    .B(_00751_),
    .C(net298),
    .ZN(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05924_ (.I(_00752_),
    .Z(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05925_ (.I(_00753_),
    .Z(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05926_ (.A1(_00749_),
    .A2(_00754_),
    .ZN(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05927_ (.I(_00755_),
    .Z(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05928_ (.A1(\as2650.regs[6][7] ),
    .A2(_00756_),
    .Z(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _05929_ (.A1(\as2650.insin[1] ),
    .A2(_00672_),
    .Z(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05930_ (.I(_00758_),
    .Z(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05931_ (.I(net43),
    .ZN(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05932_ (.A1(_00665_),
    .A2(_00668_),
    .B(net31),
    .ZN(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05933_ (.A1(_00760_),
    .A2(_00682_),
    .B(_00761_),
    .C(_00672_),
    .ZN(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05934_ (.I(_00762_),
    .Z(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05935_ (.A1(_00759_),
    .A2(_00763_),
    .ZN(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05936_ (.I(_00764_),
    .Z(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _05937_ (.A1(\as2650.regs[7][7] ),
    .A2(_00746_),
    .B(_00757_),
    .C(_00765_),
    .ZN(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _05938_ (.A1(_00759_),
    .A2(_00763_),
    .A3(_00742_),
    .A4(_00743_),
    .Z(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05939_ (.I(_00767_),
    .Z(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _05940_ (.A1(_00758_),
    .A2(_00762_),
    .A3(_00748_),
    .A4(_00753_),
    .Z(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05941_ (.I(_00769_),
    .Z(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05942_ (.I(_00593_),
    .Z(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _05943_ (.A1(\as2650.regs[5][7] ),
    .A2(_00768_),
    .B1(_00770_),
    .B2(\as2650.regs[4][7] ),
    .C(_00771_),
    .ZN(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05944_ (.A1(\as2650.regs[2][7] ),
    .A2(_00756_),
    .Z(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05945_ (.I(_00764_),
    .Z(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _05946_ (.A1(\as2650.regs[3][7] ),
    .A2(_00746_),
    .B(_00773_),
    .C(_00774_),
    .ZN(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05947_ (.I(_00767_),
    .Z(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05948_ (.I(_00609_),
    .Z(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05949_ (.I(_00777_),
    .Z(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _05950_ (.A1(\as2650.regs[1][7] ),
    .A2(_00776_),
    .B1(_00770_),
    .B2(\as2650.regs[0][7] ),
    .C(_00778_),
    .ZN(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _05951_ (.A1(_00766_),
    .A2(_00772_),
    .B1(_00775_),
    .B2(_00779_),
    .ZN(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05952_ (.I(_00780_),
    .Z(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05953_ (.I(_00755_),
    .Z(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05954_ (.A1(\as2650.regs[2][6] ),
    .A2(_00782_),
    .ZN(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05955_ (.I(_00745_),
    .Z(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05956_ (.I(_00784_),
    .Z(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05957_ (.A1(\as2650.regs[3][6] ),
    .A2(_00785_),
    .ZN(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05958_ (.I(_00764_),
    .Z(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05959_ (.I(_00787_),
    .Z(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05960_ (.A1(_00783_),
    .A2(_00786_),
    .B(_00788_),
    .ZN(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05961_ (.A1(_00759_),
    .A2(_00763_),
    .A3(net295),
    .A4(_00743_),
    .ZN(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05962_ (.I(_00790_),
    .Z(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05963_ (.A1(\as2650.regs[1][6] ),
    .A2(_00791_),
    .ZN(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05964_ (.A1(_00758_),
    .A2(net293),
    .A3(_00747_),
    .A4(net300),
    .ZN(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05965_ (.I(_00793_),
    .Z(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05966_ (.I(_00794_),
    .Z(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05967_ (.A1(\as2650.regs[0][6] ),
    .A2(_00795_),
    .ZN(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05968_ (.A1(_00611_),
    .A2(_00792_),
    .A3(_00796_),
    .ZN(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05969_ (.I(_00579_),
    .Z(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05970_ (.I(_00749_),
    .Z(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05971_ (.I(_00754_),
    .Z(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05972_ (.A1(\as2650.regs[6][6] ),
    .A2(_00799_),
    .A3(_00800_),
    .Z(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05973_ (.A1(_00759_),
    .A2(_00763_),
    .Z(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05974_ (.I(_00802_),
    .Z(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _05975_ (.A1(\as2650.regs[7][6] ),
    .A2(_00756_),
    .B(_00801_),
    .C(_00803_),
    .ZN(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05976_ (.I(_00790_),
    .Z(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05977_ (.A1(\as2650.regs[5][6] ),
    .A2(_00805_),
    .ZN(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05978_ (.A1(\as2650.regs[4][6] ),
    .A2(_00795_),
    .ZN(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _05979_ (.A1(_00798_),
    .A2(_00804_),
    .A3(_00806_),
    .A4(_00807_),
    .ZN(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05980_ (.A1(_00789_),
    .A2(_00797_),
    .B(_00808_),
    .ZN(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05981_ (.I(\as2650.regs[7][5] ),
    .ZN(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05982_ (.I(_00745_),
    .Z(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _05983_ (.A1(\as2650.regs[6][5] ),
    .A2(_00799_),
    .A3(_00800_),
    .ZN(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05984_ (.A1(_00810_),
    .A2(_00811_),
    .B(_00812_),
    .C(_00774_),
    .ZN(_00813_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05985_ (.I(\as2650.regs[5][5] ),
    .ZN(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05986_ (.I(_00769_),
    .Z(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05987_ (.I(\as2650.regs[4][5] ),
    .ZN(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _05988_ (.A1(_00814_),
    .A2(_00776_),
    .B1(_00815_),
    .B2(_00816_),
    .C(_00580_),
    .ZN(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05989_ (.I(\as2650.regs[2][5] ),
    .ZN(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05990_ (.I(_00742_),
    .Z(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05991_ (.I(_00744_),
    .Z(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _05992_ (.A1(\as2650.regs[3][5] ),
    .A2(_00819_),
    .A3(_00820_),
    .ZN(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05993_ (.A1(_00818_),
    .A2(_00782_),
    .B(_00821_),
    .C(_00774_),
    .ZN(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05994_ (.I(\as2650.regs[1][5] ),
    .ZN(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05995_ (.I(_00767_),
    .Z(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05996_ (.I(\as2650.regs[0][5] ),
    .ZN(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _05997_ (.A1(_00823_),
    .A2(_00824_),
    .B1(_00815_),
    .B2(_00825_),
    .C(_00778_),
    .ZN(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _05998_ (.A1(_00813_),
    .A2(_00817_),
    .B1(_00822_),
    .B2(_00826_),
    .ZN(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05999_ (.I(\as2650.regs[7][4] ),
    .ZN(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06000_ (.I(_00745_),
    .Z(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06001_ (.I(_00748_),
    .Z(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06002_ (.I(_00753_),
    .Z(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06003_ (.A1(\as2650.regs[6][4] ),
    .A2(_00830_),
    .A3(_00831_),
    .ZN(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _06004_ (.A1(_00828_),
    .A2(_00829_),
    .B(_00832_),
    .C(_00787_),
    .ZN(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06005_ (.I(\as2650.regs[5][4] ),
    .ZN(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06006_ (.I(_00769_),
    .Z(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _06007_ (.A1(_00834_),
    .A2(_00824_),
    .B1(_00835_),
    .B2(_00632_),
    .C(_00593_),
    .ZN(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06008_ (.I(\as2650.regs[2][4] ),
    .ZN(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06009_ (.A1(\as2650.regs[3][4] ),
    .A2(_00742_),
    .A3(_00744_),
    .ZN(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _06010_ (.A1(_00837_),
    .A2(_00755_),
    .B(_00838_),
    .C(_00764_),
    .ZN(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06011_ (.I(\as2650.regs[1][4] ),
    .ZN(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06012_ (.I(\as2650.regs[0][4] ),
    .ZN(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _06013_ (.A1(_00840_),
    .A2(_00767_),
    .B1(_00835_),
    .B2(_00841_),
    .C(_00610_),
    .ZN(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _06014_ (.A1(_00833_),
    .A2(_00836_),
    .B1(_00839_),
    .B2(_00842_),
    .ZN(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06015_ (.I(_00843_),
    .Z(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06016_ (.I(\as2650.regs[6][1] ),
    .ZN(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06017_ (.I(_00748_),
    .Z(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06018_ (.A1(_00846_),
    .A2(_00831_),
    .B(\as2650.regs[7][1] ),
    .ZN(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06019_ (.I(_00802_),
    .Z(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06020_ (.A1(_00845_),
    .A2(_00811_),
    .B(_00847_),
    .C(_00848_),
    .ZN(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06021_ (.I(\as2650.regs[5][1] ),
    .ZN(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06022_ (.I(_00793_),
    .Z(_00851_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06023_ (.I(\as2650.regs[4][1] ),
    .ZN(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06024_ (.A1(_00850_),
    .A2(_00805_),
    .B1(_00851_),
    .B2(_00852_),
    .C(_00610_),
    .ZN(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _06025_ (.I(\as2650.regs[2][1] ),
    .ZN(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06026_ (.A1(_00830_),
    .A2(_00831_),
    .B(\as2650.regs[3][1] ),
    .ZN(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06027_ (.A1(_00854_),
    .A2(_00811_),
    .B(_00855_),
    .C(_00848_),
    .ZN(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06028_ (.I(\as2650.regs[1][1] ),
    .ZN(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06029_ (.I(\as2650.regs[0][1] ),
    .ZN(_00858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06030_ (.I(\as2650.debug_psl[4] ),
    .Z(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06031_ (.A1(_00857_),
    .A2(_00805_),
    .B1(_00795_),
    .B2(_00858_),
    .C(_00859_),
    .ZN(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06032_ (.A1(_00849_),
    .A2(_00853_),
    .B1(_00856_),
    .B2(_00860_),
    .ZN(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06033_ (.I(\as2650.regs[6][0] ),
    .ZN(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06034_ (.A1(_00749_),
    .A2(_00754_),
    .B(\as2650.regs[7][0] ),
    .ZN(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06035_ (.I(_00802_),
    .Z(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06036_ (.A1(_00862_),
    .A2(_00784_),
    .B(_00863_),
    .C(_00864_),
    .ZN(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06037_ (.I(\as2650.regs[5][0] ),
    .ZN(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06038_ (.I(\as2650.regs[4][0] ),
    .ZN(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06039_ (.A1(_00866_),
    .A2(_00790_),
    .B1(net299),
    .B2(_00867_),
    .C(_00777_),
    .ZN(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _06040_ (.I(\as2650.regs[2][0] ),
    .ZN(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06041_ (.A1(_00749_),
    .A2(_00754_),
    .B(\as2650.regs[3][0] ),
    .ZN(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06042_ (.A1(_00869_),
    .A2(_00784_),
    .B(_00870_),
    .C(_00864_),
    .ZN(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06043_ (.I(\as2650.regs[1][0] ),
    .ZN(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06044_ (.I(_00790_),
    .Z(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06045_ (.I(\as2650.regs[0][0] ),
    .ZN(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06046_ (.A1(_00872_),
    .A2(_00873_),
    .B1(net299),
    .B2(_00874_),
    .C(_00859_),
    .ZN(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06047_ (.A1(_00865_),
    .A2(_00868_),
    .B1(_00871_),
    .B2(_00875_),
    .ZN(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06048_ (.I(\as2650.regs[6][3] ),
    .ZN(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06049_ (.I(_00753_),
    .Z(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06050_ (.A1(_00846_),
    .A2(_00878_),
    .B(\as2650.regs[7][3] ),
    .ZN(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06051_ (.A1(_00877_),
    .A2(_00784_),
    .B(_00879_),
    .C(_00864_),
    .ZN(_00880_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06052_ (.I(\as2650.regs[5][3] ),
    .ZN(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06053_ (.I(\as2650.regs[4][3] ),
    .ZN(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06054_ (.A1(_00881_),
    .A2(_00873_),
    .B1(net299),
    .B2(_00882_),
    .C(_00777_),
    .ZN(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06055_ (.I(\as2650.regs[2][3] ),
    .ZN(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06056_ (.A1(_00846_),
    .A2(_00878_),
    .B(\as2650.regs[3][3] ),
    .ZN(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06057_ (.A1(_00884_),
    .A2(_00829_),
    .B(_00885_),
    .C(_00864_),
    .ZN(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06058_ (.I(\as2650.regs[1][3] ),
    .ZN(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06059_ (.I(\as2650.regs[0][3] ),
    .ZN(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06060_ (.A1(_00887_),
    .A2(_00873_),
    .B1(_00851_),
    .B2(_00888_),
    .C(_00859_),
    .ZN(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06061_ (.A1(_00880_),
    .A2(_00883_),
    .B1(_00886_),
    .B2(_00889_),
    .ZN(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06062_ (.I(\as2650.regs[6][2] ),
    .ZN(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06063_ (.A1(_00846_),
    .A2(_00878_),
    .B(\as2650.regs[7][2] ),
    .ZN(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06064_ (.A1(_00891_),
    .A2(_00829_),
    .B(_00892_),
    .C(_00848_),
    .ZN(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06065_ (.I(\as2650.regs[5][2] ),
    .ZN(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06066_ (.I(\as2650.regs[4][2] ),
    .ZN(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06067_ (.A1(_00894_),
    .A2(_00873_),
    .B1(_00851_),
    .B2(_00895_),
    .C(_00777_),
    .ZN(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _06068_ (.I(\as2650.regs[2][2] ),
    .ZN(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06069_ (.A1(_00830_),
    .A2(_00831_),
    .B(\as2650.regs[3][2] ),
    .ZN(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06070_ (.A1(_00897_),
    .A2(_00811_),
    .B(_00898_),
    .C(_00848_),
    .ZN(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06071_ (.I(\as2650.regs[1][2] ),
    .ZN(_00900_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06072_ (.I(\as2650.regs[0][2] ),
    .ZN(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06073_ (.A1(_00900_),
    .A2(_00805_),
    .B1(_00851_),
    .B2(_00901_),
    .C(_00859_),
    .ZN(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06074_ (.A1(_00893_),
    .A2(_00896_),
    .B1(_00899_),
    .B2(_00902_),
    .ZN(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _06075_ (.A1(_00861_),
    .A2(_00876_),
    .A3(_00890_),
    .A4(_00903_),
    .Z(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _06076_ (.A1(_00809_),
    .A2(_00827_),
    .A3(_00844_),
    .A4(_00904_),
    .ZN(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06077_ (.A1(_00781_),
    .A2(_00905_),
    .Z(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _06078_ (.A1(_00739_),
    .A2(_00906_),
    .Z(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06079_ (.A1(\as2650.extend ),
    .A2(_00737_),
    .ZN(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06080_ (.A1(_00733_),
    .A2(_00908_),
    .ZN(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06081_ (.I(_00909_),
    .Z(_00910_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06082_ (.I(_00780_),
    .ZN(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06083_ (.I(_00756_),
    .Z(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06084_ (.A1(\as2650.regs[2][6] ),
    .A2(_00746_),
    .Z(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06085_ (.A1(\as2650.regs[3][6] ),
    .A2(_00912_),
    .B(_00913_),
    .C(_00803_),
    .ZN(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06086_ (.A1(_00611_),
    .A2(_00792_),
    .A3(_00796_),
    .Z(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _06087_ (.A1(_00590_),
    .A2(_00804_),
    .A3(_00806_),
    .A4(_00807_),
    .Z(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06088_ (.A1(_00914_),
    .A2(_00915_),
    .B(_00916_),
    .ZN(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06089_ (.A1(_00861_),
    .A2(_00876_),
    .A3(_00890_),
    .A4(_00903_),
    .ZN(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06090_ (.A1(_00827_),
    .A2(_00844_),
    .ZN(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06091_ (.A1(_00917_),
    .A2(_00918_),
    .A3(_00919_),
    .ZN(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06092_ (.A1(_00911_),
    .A2(_00920_),
    .Z(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06093_ (.A1(_00781_),
    .A2(_00910_),
    .ZN(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06094_ (.A1(_00910_),
    .A2(_00921_),
    .B(_00922_),
    .C(_00739_),
    .ZN(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _06095_ (.A1(_00730_),
    .A2(_00907_),
    .A3(_00923_),
    .Z(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _06096_ (.I(\as2650.indirect_cyc ),
    .ZN(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06097_ (.A1(_00652_),
    .A2(_00925_),
    .ZN(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06098_ (.I(_00926_),
    .Z(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06099_ (.I(_00927_),
    .Z(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06100_ (.A1(\as2650.cycle[2] ),
    .A2(\as2650.cycle[3] ),
    .Z(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06101_ (.I(_00929_),
    .Z(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06102_ (.A1(_00653_),
    .A2(_00642_),
    .ZN(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06103_ (.A1(_00929_),
    .A2(_00931_),
    .ZN(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06104_ (.I(_00932_),
    .Z(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06105_ (.I(_00646_),
    .ZN(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _06106_ (.A1(_00642_),
    .A2(_00934_),
    .A3(_00641_),
    .B(_00925_),
    .ZN(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06107_ (.A1(\as2650.relative_cyc ),
    .A2(_00930_),
    .A3(_00933_),
    .A4(_00935_),
    .ZN(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06108_ (.I(_00936_),
    .Z(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06109_ (.I(_00937_),
    .Z(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06110_ (.A1(\as2650.indirect_target[7] ),
    .A2(_00928_),
    .B1(_00938_),
    .B2(\as2650.PC[7] ),
    .ZN(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06111_ (.A1(\as2650.indirect_target[6] ),
    .A2(_00928_),
    .B1(_00938_),
    .B2(\as2650.PC[6] ),
    .ZN(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06112_ (.A1(\as2650.indirect_target[5] ),
    .A2(_00927_),
    .B1(_00937_),
    .B2(\as2650.PC[5] ),
    .ZN(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06113_ (.I(_00941_),
    .ZN(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06114_ (.A1(\as2650.indirect_target[4] ),
    .A2(_00927_),
    .ZN(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06115_ (.A1(\as2650.PC[4] ),
    .A2(_00937_),
    .ZN(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06116_ (.A1(_00943_),
    .A2(_00944_),
    .ZN(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06117_ (.I(\as2650.PC[3] ),
    .ZN(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _06118_ (.A1(\as2650.relative_cyc ),
    .A2(_00930_),
    .A3(_00932_),
    .A4(_00935_),
    .Z(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06119_ (.A1(\as2650.indirect_target[3] ),
    .A2(_00927_),
    .ZN(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06120_ (.A1(_00946_),
    .A2(_00947_),
    .B(_00948_),
    .ZN(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06121_ (.A1(\as2650.indirect_target[1] ),
    .A2(_00926_),
    .B1(_00936_),
    .B2(\as2650.PC[1] ),
    .ZN(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06122_ (.I(\as2650.PC[0] ),
    .ZN(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06123_ (.A1(\as2650.indirect_target[0] ),
    .A2(_00926_),
    .ZN(_00952_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06124_ (.I0(_00951_),
    .I1(_00952_),
    .S(_00947_),
    .Z(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06125_ (.I(\as2650.relative_cyc ),
    .Z(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06126_ (.I(_00935_),
    .Z(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06127_ (.A1(_00954_),
    .A2(_00955_),
    .Z(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06128_ (.A1(_00653_),
    .A2(_00644_),
    .A3(_00930_),
    .ZN(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06129_ (.A1(_00956_),
    .A2(_00957_),
    .ZN(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06130_ (.A1(\as2650.indirect_target[2] ),
    .A2(_00926_),
    .B1(_00937_),
    .B2(\as2650.PC[2] ),
    .ZN(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06131_ (.A1(_00950_),
    .A2(_00953_),
    .A3(_00958_),
    .A4(_00959_),
    .ZN(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06132_ (.A1(_00942_),
    .A2(_00945_),
    .A3(_00949_),
    .A4(_00960_),
    .ZN(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06133_ (.A1(_00940_),
    .A2(_00961_),
    .Z(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06134_ (.A1(_00939_),
    .A2(_00962_),
    .ZN(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06135_ (.I(_00657_),
    .Z(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06136_ (.A1(_00939_),
    .A2(_00962_),
    .ZN(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06137_ (.A1(_00964_),
    .A2(_00965_),
    .ZN(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06138_ (.I(_00933_),
    .Z(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06139_ (.A1(\as2650.instruction_args_latch[7] ),
    .A2(_00967_),
    .ZN(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06140_ (.A1(_00963_),
    .A2(_00966_),
    .B(_00968_),
    .ZN(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _06141_ (.A1(_00924_),
    .A2(_00969_),
    .ZN(_00970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06142_ (.A1(_00660_),
    .A2(_00728_),
    .ZN(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06143_ (.I(_00971_),
    .Z(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06144_ (.I(_00876_),
    .Z(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06145_ (.I(_00890_),
    .Z(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06146_ (.A1(_00861_),
    .A2(_00973_),
    .A3(_00974_),
    .A4(_00903_),
    .Z(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06147_ (.I(_00827_),
    .Z(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06148_ (.I(_00843_),
    .Z(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06149_ (.A1(_00976_),
    .A2(_00977_),
    .Z(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06150_ (.A1(_00975_),
    .A2(_00978_),
    .B(_00809_),
    .ZN(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06151_ (.I(_00909_),
    .Z(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06152_ (.I(_00809_),
    .Z(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06153_ (.A1(_00980_),
    .A2(_00981_),
    .ZN(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06154_ (.A1(_00910_),
    .A2(_00920_),
    .A3(_00979_),
    .B(_00982_),
    .ZN(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _06155_ (.A1(_00827_),
    .A2(_00844_),
    .A3(_00904_),
    .Z(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06156_ (.A1(_00917_),
    .A2(_00984_),
    .Z(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _06157_ (.A1(_00734_),
    .A2(_00737_),
    .Z(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06158_ (.I(_00986_),
    .Z(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _06159_ (.I0(_00983_),
    .I1(_00985_),
    .S(_00987_),
    .Z(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06160_ (.A1(_00972_),
    .A2(_00988_),
    .ZN(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06161_ (.I(_00933_),
    .Z(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06162_ (.A1(_00940_),
    .A2(_00961_),
    .ZN(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06163_ (.A1(\as2650.instruction_args_latch[6] ),
    .A2(_00967_),
    .ZN(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06164_ (.A1(_00990_),
    .A2(_00991_),
    .B(_00992_),
    .ZN(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06165_ (.I(_00993_),
    .ZN(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06166_ (.A1(_00989_),
    .A2(_00994_),
    .Z(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06167_ (.A1(_00862_),
    .A2(_00799_),
    .A3(_00800_),
    .ZN(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06168_ (.A1(\as2650.regs[7][0] ),
    .A2(_00746_),
    .B(_00996_),
    .C(_00765_),
    .ZN(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _06169_ (.A1(\as2650.regs[5][0] ),
    .A2(_00768_),
    .B1(_00770_),
    .B2(\as2650.regs[4][0] ),
    .C(_00580_),
    .ZN(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06170_ (.I(\as2650.regs[3][0] ),
    .ZN(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06171_ (.A1(_00999_),
    .A2(_00819_),
    .A3(_00820_),
    .ZN(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06172_ (.A1(\as2650.regs[2][0] ),
    .A2(_00782_),
    .B(_01000_),
    .C(_00774_),
    .ZN(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06173_ (.I(\as2650.regs[0][0] ),
    .Z(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _06174_ (.A1(\as2650.regs[1][0] ),
    .A2(_00776_),
    .B1(_00815_),
    .B2(_01002_),
    .C(_00778_),
    .ZN(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _06175_ (.A1(_00997_),
    .A2(_00998_),
    .B1(_01001_),
    .B2(_01003_),
    .ZN(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06176_ (.I(_01004_),
    .Z(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06177_ (.A1(_00738_),
    .A2(_00909_),
    .ZN(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06178_ (.A1(_01005_),
    .A2(_01006_),
    .Z(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _06179_ (.I(\as2650.instruction_args_latch[0] ),
    .ZN(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06180_ (.A1(_00953_),
    .A2(_00958_),
    .Z(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06181_ (.A1(_00953_),
    .A2(_00958_),
    .Z(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06182_ (.A1(_00657_),
    .A2(_01010_),
    .ZN(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _06183_ (.A1(_01008_),
    .A2(_00657_),
    .B1(_01009_),
    .B2(_01011_),
    .ZN(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06184_ (.A1(_00730_),
    .A2(_01007_),
    .A3(_01012_),
    .Z(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06185_ (.A1(_00845_),
    .A2(_00830_),
    .A3(_00878_),
    .ZN(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06186_ (.A1(\as2650.regs[7][1] ),
    .A2(_00829_),
    .B(_01014_),
    .C(_00787_),
    .ZN(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _06187_ (.A1(\as2650.regs[5][1] ),
    .A2(_00824_),
    .B1(_00815_),
    .B2(\as2650.regs[4][1] ),
    .C(_00593_),
    .ZN(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06188_ (.I(\as2650.regs[3][1] ),
    .ZN(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06189_ (.A1(_01017_),
    .A2(_00819_),
    .A3(_00744_),
    .ZN(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06190_ (.A1(\as2650.regs[2][1] ),
    .A2(_00755_),
    .B(_01018_),
    .C(_00787_),
    .ZN(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06191_ (.I(\as2650.regs[0][1] ),
    .Z(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _06192_ (.A1(\as2650.regs[1][1] ),
    .A2(_00824_),
    .B1(_00835_),
    .B2(_01020_),
    .C(_00610_),
    .ZN(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _06193_ (.A1(_01015_),
    .A2(_01016_),
    .B1(_01019_),
    .B2(_01021_),
    .ZN(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06194_ (.I(_01022_),
    .Z(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06195_ (.A1(_01023_),
    .A2(_00876_),
    .Z(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _06196_ (.A1(_00733_),
    .A2(_00908_),
    .Z(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06197_ (.A1(_01025_),
    .A2(_01005_),
    .B(_00738_),
    .ZN(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06198_ (.A1(_01024_),
    .A2(_01026_),
    .ZN(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _06199_ (.A1(_00950_),
    .A2(_01010_),
    .ZN(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06200_ (.I(_00933_),
    .Z(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06201_ (.A1(\as2650.instruction_args_latch[1] ),
    .A2(_01029_),
    .ZN(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _06202_ (.A1(_00972_),
    .A2(_01027_),
    .B1(_01028_),
    .B2(_00990_),
    .C(_01030_),
    .ZN(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06203_ (.A1(_01024_),
    .A2(_01026_),
    .Z(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06204_ (.A1(_01029_),
    .A2(_01028_),
    .B(_01030_),
    .ZN(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _06205_ (.A1(_00730_),
    .A2(_01032_),
    .A3(_01033_),
    .Z(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06206_ (.A1(_01013_),
    .A2(_01031_),
    .B(_01034_),
    .ZN(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06207_ (.A1(_00891_),
    .A2(_00799_),
    .A3(_00800_),
    .ZN(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06208_ (.A1(\as2650.regs[7][2] ),
    .A2(_00785_),
    .B(_01036_),
    .C(_00765_),
    .ZN(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06209_ (.I(_00835_),
    .Z(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _06210_ (.A1(\as2650.regs[5][2] ),
    .A2(_00768_),
    .B1(_01038_),
    .B2(\as2650.regs[4][2] ),
    .C(_00771_),
    .ZN(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06211_ (.I(\as2650.regs[3][2] ),
    .ZN(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06212_ (.A1(_01040_),
    .A2(_00819_),
    .A3(_00820_),
    .ZN(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06213_ (.A1(\as2650.regs[2][2] ),
    .A2(_00782_),
    .B(_01041_),
    .C(_00765_),
    .ZN(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06214_ (.I(\as2650.regs[0][2] ),
    .Z(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _06215_ (.A1(\as2650.regs[1][2] ),
    .A2(_00776_),
    .B1(_00770_),
    .B2(_01043_),
    .C(_00778_),
    .ZN(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _06216_ (.A1(_01037_),
    .A2(_01039_),
    .B1(_01042_),
    .B2(_01044_),
    .ZN(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06217_ (.A1(_01022_),
    .A2(_01004_),
    .A3(_01045_),
    .ZN(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06218_ (.I(_01046_),
    .Z(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06219_ (.I(_00861_),
    .Z(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06220_ (.I(_00903_),
    .Z(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06221_ (.A1(_01048_),
    .A2(_00973_),
    .B(_01049_),
    .ZN(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06222_ (.A1(_00909_),
    .A2(_01049_),
    .ZN(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _06223_ (.A1(_00980_),
    .A2(_01047_),
    .A3(_01050_),
    .B(_01051_),
    .ZN(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06224_ (.A1(_01022_),
    .A2(_01004_),
    .A3(_01045_),
    .ZN(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06225_ (.A1(_01048_),
    .A2(_00973_),
    .B(_01049_),
    .ZN(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06226_ (.I(_00738_),
    .Z(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06227_ (.A1(_01053_),
    .A2(_01054_),
    .B(_01055_),
    .ZN(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06228_ (.A1(_00739_),
    .A2(_01052_),
    .B(_01056_),
    .C(_00971_),
    .ZN(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06229_ (.A1(_00950_),
    .A2(_01010_),
    .ZN(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06230_ (.A1(_01058_),
    .A2(_00959_),
    .Z(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06231_ (.A1(\as2650.instruction_args_latch[2] ),
    .A2(_01029_),
    .ZN(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06232_ (.A1(_00967_),
    .A2(_01059_),
    .B(_01060_),
    .ZN(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06233_ (.I(_01061_),
    .Z(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06234_ (.A1(_01057_),
    .A2(_01062_),
    .ZN(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06235_ (.I(_01057_),
    .Z(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06236_ (.A1(_01064_),
    .A2(_01061_),
    .ZN(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06237_ (.A1(_01035_),
    .A2(_01063_),
    .B(_01065_),
    .ZN(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06238_ (.I(_00918_),
    .Z(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06239_ (.A1(_00974_),
    .A2(_01046_),
    .B(_01067_),
    .C(_01025_),
    .ZN(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06240_ (.A1(_00980_),
    .A2(_00974_),
    .ZN(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _06241_ (.A1(_01055_),
    .A2(_01068_),
    .A3(_01069_),
    .Z(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06242_ (.A1(_00880_),
    .A2(_00883_),
    .ZN(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06243_ (.A1(_00886_),
    .A2(_00889_),
    .ZN(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06244_ (.A1(_01071_),
    .A2(_01072_),
    .ZN(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06245_ (.A1(_01073_),
    .A2(_01053_),
    .Z(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06246_ (.A1(_01055_),
    .A2(_01074_),
    .ZN(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06247_ (.A1(_01070_),
    .A2(_01075_),
    .B(_00729_),
    .ZN(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06248_ (.A1(_00949_),
    .A2(_00960_),
    .Z(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06249_ (.A1(_00949_),
    .A2(_00960_),
    .ZN(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06250_ (.A1(_01029_),
    .A2(_01077_),
    .A3(_01078_),
    .ZN(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06251_ (.A1(\as2650.instruction_args_latch[3] ),
    .A2(_00990_),
    .B(_01079_),
    .ZN(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06252_ (.A1(_01076_),
    .A2(_01080_),
    .Z(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06253_ (.A1(_01076_),
    .A2(_01080_),
    .ZN(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06254_ (.A1(_01066_),
    .A2(_01081_),
    .B(_01082_),
    .ZN(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06255_ (.A1(_01067_),
    .A2(_00919_),
    .ZN(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06256_ (.A1(_00975_),
    .A2(_00977_),
    .B(_00976_),
    .ZN(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06257_ (.I(_00976_),
    .Z(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06258_ (.A1(_00980_),
    .A2(_01086_),
    .ZN(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _06259_ (.A1(_00910_),
    .A2(_01084_),
    .A3(_01085_),
    .B(_01087_),
    .ZN(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06260_ (.I(_00844_),
    .Z(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06261_ (.A1(_01089_),
    .A2(_00904_),
    .B(_00976_),
    .ZN(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06262_ (.A1(_00984_),
    .A2(_01090_),
    .B(_01055_),
    .ZN(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06263_ (.A1(_00739_),
    .A2(_01088_),
    .B(_01091_),
    .C(_00971_),
    .ZN(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06264_ (.A1(_00945_),
    .A2(_01077_),
    .B(_00942_),
    .ZN(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06265_ (.A1(_00964_),
    .A2(_00961_),
    .ZN(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06266_ (.A1(\as2650.instruction_args_latch[5] ),
    .A2(_00967_),
    .ZN(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06267_ (.A1(_01093_),
    .A2(_01094_),
    .B(_01095_),
    .ZN(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06268_ (.A1(_01092_),
    .A2(_01096_),
    .Z(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _06269_ (.A1(_00977_),
    .A2(_00904_),
    .ZN(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06270_ (.A1(_01067_),
    .A2(_00977_),
    .Z(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06271_ (.A1(_01025_),
    .A2(_01089_),
    .ZN(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06272_ (.A1(_01025_),
    .A2(_01099_),
    .B(_01100_),
    .C(_00986_),
    .ZN(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06273_ (.A1(_00987_),
    .A2(_01098_),
    .B(_01101_),
    .C(_00972_),
    .ZN(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06274_ (.A1(_00945_),
    .A2(_01077_),
    .Z(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06275_ (.I0(\as2650.instruction_args_latch[4] ),
    .I1(_01103_),
    .S(_00964_),
    .Z(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06276_ (.A1(_01104_),
    .A2(_01102_),
    .Z(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06277_ (.A1(_01105_),
    .A2(_01097_),
    .ZN(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06278_ (.A1(_00970_),
    .A2(_00995_),
    .A3(_01083_),
    .A4(_01106_),
    .ZN(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06279_ (.I(_01107_),
    .Z(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06280_ (.A1(_01092_),
    .A2(_01096_),
    .Z(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06281_ (.A1(_01102_),
    .A2(_01104_),
    .Z(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06282_ (.A1(_01092_),
    .A2(_01096_),
    .Z(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06283_ (.A1(_01109_),
    .A2(_01110_),
    .B(_01111_),
    .ZN(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06284_ (.A1(_00972_),
    .A2(_00988_),
    .A3(_00994_),
    .ZN(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06285_ (.A1(_00924_),
    .A2(_00969_),
    .B(_01113_),
    .ZN(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06286_ (.A1(_00924_),
    .A2(_00969_),
    .ZN(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _06287_ (.A1(_00970_),
    .A2(_00995_),
    .A3(_01112_),
    .B1(_01114_),
    .B2(_01115_),
    .ZN(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06288_ (.I(_01116_),
    .Z(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06289_ (.I(_00990_),
    .Z(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06290_ (.I(_01118_),
    .Z(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06291_ (.A1(\as2650.indirect_target[8] ),
    .A2(_00928_),
    .B1(_00938_),
    .B2(\as2650.PC[8] ),
    .ZN(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06292_ (.A1(_00939_),
    .A2(_00940_),
    .A3(_00961_),
    .A4(_01120_),
    .ZN(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06293_ (.I(_00928_),
    .Z(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06294_ (.A1(\as2650.indirect_target[9] ),
    .A2(_01122_),
    .ZN(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06295_ (.I(_00938_),
    .Z(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06296_ (.A1(\as2650.PC[9] ),
    .A2(_01124_),
    .ZN(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06297_ (.A1(_01123_),
    .A2(_01125_),
    .ZN(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06298_ (.A1(_01121_),
    .A2(_01126_),
    .ZN(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06299_ (.I(_01127_),
    .Z(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06300_ (.A1(\as2650.indirect_target[10] ),
    .A2(_01122_),
    .B1(_01124_),
    .B2(\as2650.PC[10] ),
    .ZN(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06301_ (.I(_01129_),
    .Z(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06302_ (.A1(\as2650.indirect_target[11] ),
    .A2(_01122_),
    .B1(_01124_),
    .B2(\as2650.PC[11] ),
    .ZN(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06303_ (.A1(_01128_),
    .A2(_01130_),
    .B(_01131_),
    .ZN(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06304_ (.I(_01118_),
    .Z(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06305_ (.A1(_01127_),
    .A2(_01130_),
    .A3(_01131_),
    .ZN(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06306_ (.A1(_01133_),
    .A2(_01134_),
    .ZN(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06307_ (.A1(\as2650.instruction_args_latch[11] ),
    .A2(_01119_),
    .B1(_01132_),
    .B2(_01135_),
    .ZN(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06308_ (.A1(_01128_),
    .A2(_01130_),
    .ZN(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06309_ (.A1(_01128_),
    .A2(_01130_),
    .Z(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06310_ (.A1(\as2650.instruction_args_latch[10] ),
    .A2(_01118_),
    .ZN(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06311_ (.A1(_01133_),
    .A2(_01137_),
    .A3(_01138_),
    .B(_01139_),
    .ZN(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06312_ (.A1(_00963_),
    .A2(_01120_),
    .Z(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06313_ (.A1(\as2650.instruction_args_latch[8] ),
    .A2(_01118_),
    .ZN(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06314_ (.A1(_01133_),
    .A2(_01141_),
    .B(_01142_),
    .ZN(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06315_ (.I(\as2650.instruction_args_latch[9] ),
    .ZN(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06316_ (.I(_00964_),
    .Z(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06317_ (.A1(_01121_),
    .A2(_01126_),
    .ZN(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06318_ (.A1(_01145_),
    .A2(_01128_),
    .ZN(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _06319_ (.A1(_01144_),
    .A2(_01145_),
    .B1(_01146_),
    .B2(_01147_),
    .ZN(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06320_ (.A1(_01140_),
    .A2(_01143_),
    .A3(_01148_),
    .ZN(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06321_ (.A1(_01136_),
    .A2(_01149_),
    .ZN(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06322_ (.A1(_01108_),
    .A2(_01117_),
    .B(_01150_),
    .ZN(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06323_ (.I(_01122_),
    .Z(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06324_ (.I(_01124_),
    .Z(_01153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06325_ (.A1(\as2650.indirect_target[12] ),
    .A2(_01152_),
    .B1(_01153_),
    .B2(\as2650.PC[12] ),
    .ZN(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06326_ (.A1(_01134_),
    .A2(_01154_),
    .Z(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06327_ (.A1(\as2650.instruction_args_latch[12] ),
    .A2(_01133_),
    .ZN(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06328_ (.A1(_01119_),
    .A2(_01155_),
    .B(_01156_),
    .ZN(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06329_ (.A1(_01151_),
    .A2(_01157_),
    .Z(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06330_ (.I(_00649_),
    .Z(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06331_ (.I(_01159_),
    .Z(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06332_ (.A1(\as2650.ivectors_base[8] ),
    .A2(_01160_),
    .ZN(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06333_ (.A1(_00651_),
    .A2(_01158_),
    .B(_01161_),
    .ZN(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06334_ (.A1(\as2650.last_addr[12] ),
    .A2(_01162_),
    .Z(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06335_ (.I(_01145_),
    .Z(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06336_ (.A1(_01127_),
    .A2(_01129_),
    .A3(_01131_),
    .A4(_01154_),
    .ZN(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06337_ (.A1(\as2650.indirect_target[13] ),
    .A2(_01152_),
    .B1(_01153_),
    .B2(\as2650.page_reg[0] ),
    .ZN(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06338_ (.A1(_01165_),
    .A2(_01166_),
    .Z(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06339_ (.A1(_00658_),
    .A2(_00708_),
    .ZN(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06340_ (.I(_01168_),
    .Z(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06341_ (.A1(_00735_),
    .A2(_01168_),
    .ZN(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06342_ (.A1(\as2650.page_reg[0] ),
    .A2(_01169_),
    .B(_01170_),
    .C(_01145_),
    .ZN(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06343_ (.A1(_01164_),
    .A2(_01167_),
    .B(_01171_),
    .ZN(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06344_ (.I(_01172_),
    .ZN(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06345_ (.A1(_01108_),
    .A2(_01117_),
    .B(_01150_),
    .C(_01157_),
    .ZN(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06346_ (.A1(_01173_),
    .A2(_01174_),
    .Z(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06347_ (.A1(_00643_),
    .A2(_00934_),
    .ZN(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06348_ (.A1(_00640_),
    .A2(_01176_),
    .ZN(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06349_ (.I(_01177_),
    .Z(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06350_ (.I(_01178_),
    .Z(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06351_ (.A1(_01157_),
    .A2(_01172_),
    .Z(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06352_ (.A1(_01107_),
    .A2(_01116_),
    .B(_01150_),
    .C(_01180_),
    .ZN(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06353_ (.A1(_01179_),
    .A2(_01181_),
    .ZN(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06354_ (.A1(\as2650.ivectors_base[9] ),
    .A2(_01160_),
    .ZN(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06355_ (.A1(_01175_),
    .A2(_01182_),
    .B(_01183_),
    .ZN(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06356_ (.A1(\as2650.last_addr[13] ),
    .A2(_01184_),
    .Z(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06357_ (.A1(_01163_),
    .A2(_01185_),
    .ZN(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06358_ (.I(_01119_),
    .Z(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06359_ (.A1(_01187_),
    .A2(_01137_),
    .A3(_01138_),
    .Z(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06360_ (.A1(_01108_),
    .A2(_01117_),
    .B(_01143_),
    .C(_01148_),
    .ZN(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06361_ (.A1(_01139_),
    .A2(_01188_),
    .A3(_01189_),
    .Z(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06362_ (.I(_01177_),
    .Z(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06363_ (.I(_01149_),
    .ZN(_01192_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06364_ (.A1(_01107_),
    .A2(_01117_),
    .B(_01192_),
    .ZN(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06365_ (.A1(_01191_),
    .A2(_01193_),
    .ZN(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06366_ (.I(_00649_),
    .Z(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06367_ (.A1(\as2650.ivectors_base[6] ),
    .A2(_01195_),
    .ZN(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06368_ (.A1(_01190_),
    .A2(_01194_),
    .B(_01196_),
    .ZN(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06369_ (.A1(\as2650.last_addr[10] ),
    .A2(_01197_),
    .Z(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06370_ (.A1(_01136_),
    .A2(_01193_),
    .ZN(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06371_ (.A1(\as2650.ivectors_base[7] ),
    .A2(_01195_),
    .ZN(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06372_ (.A1(_01160_),
    .A2(_01199_),
    .B(_01200_),
    .ZN(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06373_ (.A1(\as2650.last_addr[11] ),
    .A2(_01201_),
    .Z(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _06374_ (.A1(_01108_),
    .A2(_01116_),
    .Z(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06375_ (.A1(_01203_),
    .A2(_01143_),
    .B(_01148_),
    .ZN(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06376_ (.A1(_01191_),
    .A2(_01189_),
    .ZN(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06377_ (.A1(\as2650.ivectors_base[5] ),
    .A2(_00650_),
    .ZN(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06378_ (.A1(_01204_),
    .A2(_01205_),
    .B(_01206_),
    .ZN(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06379_ (.A1(\as2650.last_addr[9] ),
    .A2(_01207_),
    .Z(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06380_ (.A1(_01203_),
    .A2(_01143_),
    .ZN(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06381_ (.A1(\as2650.ivectors_base[4] ),
    .A2(_01195_),
    .ZN(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06382_ (.A1(_01160_),
    .A2(_01209_),
    .B(_01210_),
    .ZN(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06383_ (.A1(_01211_),
    .A2(\as2650.last_addr[8] ),
    .Z(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06384_ (.A1(_01198_),
    .A2(_01202_),
    .A3(_01208_),
    .A4(_01212_),
    .ZN(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06385_ (.A1(\as2650.ivectors_base[11] ),
    .A2(_00651_),
    .Z(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06386_ (.A1(\as2650.page_reg[1] ),
    .A2(_01169_),
    .ZN(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06387_ (.A1(_00731_),
    .A2(_01169_),
    .B(_01215_),
    .ZN(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06388_ (.I(_01166_),
    .ZN(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06389_ (.A1(_01165_),
    .A2(_01217_),
    .ZN(_01218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06390_ (.A1(\as2650.indirect_target[14] ),
    .A2(_01152_),
    .B1(_01153_),
    .B2(\as2650.page_reg[1] ),
    .ZN(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06391_ (.A1(_01218_),
    .A2(_01219_),
    .ZN(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06392_ (.A1(_01218_),
    .A2(_01219_),
    .ZN(_01221_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06393_ (.A1(_01187_),
    .A2(_01221_),
    .ZN(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06394_ (.A1(_01187_),
    .A2(_01216_),
    .B1(_01220_),
    .B2(_01222_),
    .ZN(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06395_ (.I(_01164_),
    .Z(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06396_ (.I(_01153_),
    .Z(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06397_ (.A1(\as2650.indirect_target[15] ),
    .A2(_01152_),
    .B1(_01225_),
    .B2(\as2650.page_reg[2] ),
    .ZN(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06398_ (.A1(_01221_),
    .A2(_01226_),
    .Z(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06399_ (.I(_01169_),
    .Z(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06400_ (.I0(\as2650.instruction_args_latch[15] ),
    .I1(\as2650.page_reg[2] ),
    .S(_01228_),
    .Z(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06401_ (.A1(_01164_),
    .A2(_01229_),
    .ZN(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06402_ (.A1(_01224_),
    .A2(_01227_),
    .B(_01230_),
    .ZN(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06403_ (.A1(_01181_),
    .A2(_01223_),
    .A3(_01231_),
    .Z(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06404_ (.A1(_01181_),
    .A2(_01223_),
    .B(_01231_),
    .ZN(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06405_ (.A1(_01232_),
    .A2(_01233_),
    .B(_00651_),
    .ZN(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06406_ (.A1(_01214_),
    .A2(_01234_),
    .B(\as2650.last_addr[15] ),
    .ZN(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06407_ (.A1(\as2650.last_addr[15] ),
    .A2(_01214_),
    .A3(_01234_),
    .Z(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06408_ (.A1(_01181_),
    .A2(_01223_),
    .Z(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06409_ (.A1(\as2650.ivectors_base[10] ),
    .A2(_01159_),
    .Z(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06410_ (.A1(_01179_),
    .A2(_01237_),
    .B(_01238_),
    .ZN(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06411_ (.A1(\as2650.last_addr[14] ),
    .A2(_01239_),
    .ZN(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06412_ (.A1(_01235_),
    .A2(_01236_),
    .B(_01240_),
    .ZN(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06413_ (.A1(_01186_),
    .A2(_01213_),
    .A3(_01241_),
    .Z(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06414_ (.I(_00655_),
    .Z(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06415_ (.I(_00641_),
    .Z(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06416_ (.A1(_01244_),
    .A2(_01176_),
    .ZN(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06417_ (.A1(_01243_),
    .A2(_00956_),
    .B(_01245_),
    .ZN(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06418_ (.A1(_01242_),
    .A2(_01246_),
    .Z(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06419_ (.I(_01247_),
    .ZN(_01248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06420_ (.I(_01248_),
    .Z(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06421_ (.I(_01249_),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06422_ (.A1(wb_reset_override),
    .A2(wb_reset_override_en),
    .ZN(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06423_ (.A1(wb_reset_override_en),
    .A2(net25),
    .B(_01250_),
    .ZN(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06424_ (.A1(net50),
    .A2(_01251_),
    .ZN(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _06425_ (.I(_01252_),
    .ZN(net206));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06426_ (.I(_00730_),
    .Z(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06427_ (.I(_01007_),
    .Z(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06428_ (.A1(_01253_),
    .A2(_01254_),
    .A3(_01012_),
    .ZN(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06429_ (.I(_01032_),
    .Z(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06430_ (.A1(_01253_),
    .A2(_01256_),
    .B(_01033_),
    .ZN(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06431_ (.A1(_01253_),
    .A2(_01256_),
    .A3(_01033_),
    .ZN(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06432_ (.A1(_01255_),
    .A2(_01257_),
    .B(_01258_),
    .ZN(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06433_ (.A1(_01064_),
    .A2(_01062_),
    .A3(_01259_),
    .Z(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06434_ (.A1(\as2650.irqs_latch[6] ),
    .A2(\as2650.irqs_latch[7] ),
    .A3(_01178_),
    .ZN(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06435_ (.A1(\as2650.irqs_latch[4] ),
    .A2(\as2650.irqs_latch[5] ),
    .ZN(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06436_ (.A1(\as2650.irqs_latch[2] ),
    .A2(\as2650.irqs_latch[3] ),
    .B(_01262_),
    .ZN(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06437_ (.A1(_01261_),
    .A2(_01263_),
    .ZN(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06438_ (.A1(_00650_),
    .A2(_01260_),
    .B(_01264_),
    .ZN(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06439_ (.A1(_01253_),
    .A2(_01254_),
    .B(_01012_),
    .ZN(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06440_ (.A1(_01013_),
    .A2(_01266_),
    .Z(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06441_ (.A1(_00654_),
    .A2(_01177_),
    .ZN(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06442_ (.A1(_01178_),
    .A2(_01267_),
    .B(_01268_),
    .ZN(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06443_ (.A1(\as2650.last_addr[0] ),
    .A2(_01269_),
    .Z(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06444_ (.A1(_01258_),
    .A2(_01031_),
    .B(_01013_),
    .ZN(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _06445_ (.A1(_01034_),
    .A2(_01255_),
    .A3(_01257_),
    .B(_01177_),
    .ZN(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06446_ (.I(\as2650.irqs_latch[2] ),
    .ZN(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06447_ (.A1(\as2650.irqs_latch[1] ),
    .A2(_01273_),
    .B(\as2650.irqs_latch[3] ),
    .ZN(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06448_ (.A1(\as2650.irqs_latch[4] ),
    .A2(_01274_),
    .ZN(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06449_ (.A1(\as2650.irqs_latch[5] ),
    .A2(_01275_),
    .ZN(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06450_ (.A1(\as2650.irqs_latch[6] ),
    .A2(_01276_),
    .ZN(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06451_ (.A1(\as2650.irqs_latch[7] ),
    .A2(_01277_),
    .B(_00648_),
    .ZN(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06452_ (.A1(_01271_),
    .A2(_01272_),
    .B(_01278_),
    .ZN(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06453_ (.A1(\as2650.last_addr[1] ),
    .A2(_01279_),
    .Z(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06454_ (.A1(\as2650.last_addr[2] ),
    .A2(_01265_),
    .B(_01270_),
    .C(_01280_),
    .ZN(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06455_ (.A1(\as2650.last_addr[2] ),
    .A2(_01265_),
    .B(_01281_),
    .ZN(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06456_ (.A1(_01064_),
    .A2(_01062_),
    .Z(_01283_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06457_ (.A1(_01064_),
    .A2(_01062_),
    .Z(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06458_ (.A1(_01259_),
    .A2(_01283_),
    .B(_01284_),
    .ZN(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06459_ (.A1(_01285_),
    .A2(_01081_),
    .Z(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06460_ (.A1(_01261_),
    .A2(_01262_),
    .B1(_01286_),
    .B2(_01191_),
    .ZN(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06461_ (.A1(\as2650.last_addr[3] ),
    .A2(_01287_),
    .Z(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06462_ (.A1(_01076_),
    .A2(_01080_),
    .Z(_01289_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06463_ (.A1(_01076_),
    .A2(_01080_),
    .Z(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06464_ (.A1(_01285_),
    .A2(_01289_),
    .B(_01290_),
    .ZN(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06465_ (.A1(_01291_),
    .A2(_01105_),
    .Z(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06466_ (.A1(_01291_),
    .A2(_01105_),
    .B(_01178_),
    .ZN(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06467_ (.A1(\as2650.ivectors_base[0] ),
    .A2(_01159_),
    .ZN(_01294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06468_ (.A1(_01292_),
    .A2(_01293_),
    .B(_01294_),
    .ZN(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06469_ (.A1(\as2650.last_addr[4] ),
    .A2(_01295_),
    .Z(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06470_ (.A1(_01282_),
    .A2(_01288_),
    .A3(_01296_),
    .ZN(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06471_ (.I(\as2650.ivectors_base[1] ),
    .ZN(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06472_ (.A1(_01110_),
    .A2(_01292_),
    .ZN(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06473_ (.A1(_01097_),
    .A2(_01299_),
    .Z(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06474_ (.I0(_01298_),
    .I1(_01300_),
    .S(_01191_),
    .Z(_01301_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06475_ (.A1(\as2650.last_addr[5] ),
    .A2(_01301_),
    .Z(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06476_ (.A1(\as2650.ivectors_base[2] ),
    .A2(_01159_),
    .ZN(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06477_ (.A1(_00989_),
    .A2(_00993_),
    .Z(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06478_ (.A1(_01083_),
    .A2(_01106_),
    .B(_01112_),
    .ZN(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06479_ (.A1(_01304_),
    .A2(_01305_),
    .B(_00649_),
    .ZN(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06480_ (.A1(_01304_),
    .A2(_01305_),
    .B(_01306_),
    .ZN(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06481_ (.A1(_01303_),
    .A2(_01307_),
    .ZN(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06482_ (.A1(\as2650.last_addr[6] ),
    .A2(_01308_),
    .ZN(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06483_ (.A1(_01304_),
    .A2(_01305_),
    .B(_01113_),
    .ZN(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06484_ (.A1(net301),
    .A2(_01310_),
    .ZN(_01311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06485_ (.A1(\as2650.ivectors_base[3] ),
    .A2(_00650_),
    .ZN(_01312_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06486_ (.A1(_01195_),
    .A2(_01311_),
    .B(_01312_),
    .ZN(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06487_ (.A1(\as2650.last_addr[7] ),
    .A2(_01313_),
    .ZN(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _06488_ (.A1(_01297_),
    .A2(_01302_),
    .A3(_01309_),
    .A4(_01314_),
    .Z(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06489_ (.A1(_01246_),
    .A2(_01315_),
    .ZN(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06490_ (.A1(_01242_),
    .A2(_01316_),
    .ZN(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06491_ (.I(_01317_),
    .ZN(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06492_ (.I(_01318_),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06493_ (.A1(_00771_),
    .A2(_00867_),
    .ZN(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06494_ (.A1(_00798_),
    .A2(_01002_),
    .B(_01319_),
    .ZN(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06495_ (.I(_01320_),
    .ZN(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06496_ (.I(_01321_),
    .Z(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06497_ (.I(_01322_),
    .Z(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06498_ (.I(_01323_),
    .Z(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06499_ (.I(_01324_),
    .Z(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06500_ (.I(_01325_),
    .Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06501_ (.I0(_01020_),
    .I1(\as2650.regs[4][1] ),
    .S(_00581_),
    .Z(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06502_ (.I(_01326_),
    .Z(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06503_ (.I(_01327_),
    .Z(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06504_ (.I(_01328_),
    .Z(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06505_ (.I(_01329_),
    .Z(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06506_ (.I(_01330_),
    .Z(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06507_ (.I(_01331_),
    .Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06508_ (.A1(_00771_),
    .A2(_00895_),
    .ZN(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06509_ (.A1(_00798_),
    .A2(_01043_),
    .B(_01332_),
    .ZN(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06510_ (.I(_01333_),
    .ZN(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06511_ (.I(_01334_),
    .Z(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06512_ (.I(_01335_),
    .Z(_01336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06513_ (.I(_01336_),
    .Z(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06514_ (.I(_01337_),
    .Z(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06515_ (.I(_01338_),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06516_ (.I0(\as2650.regs[0][3] ),
    .I1(\as2650.regs[4][3] ),
    .S(_00798_),
    .Z(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06517_ (.I(_01339_),
    .Z(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06518_ (.I(_01340_),
    .Z(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06519_ (.I(_01341_),
    .Z(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06520_ (.I(_01342_),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _06521_ (.I(wb_io3_test),
    .ZN(net148));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06522_ (.A1(_01186_),
    .A2(net294),
    .A3(_01241_),
    .A4(_01315_),
    .ZN(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06523_ (.I(_01343_),
    .Z(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06524_ (.I(_01344_),
    .Z(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06525_ (.I(_01345_),
    .Z(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06526_ (.I(_01346_),
    .Z(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06527_ (.I(_01347_),
    .Z(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06528_ (.A1(\as2650.warmup[0] ),
    .A2(\as2650.warmup[1] ),
    .A3(net206),
    .Z(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06529_ (.I(_01349_),
    .Z(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06530_ (.I(_01350_),
    .Z(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06531_ (.I(_01351_),
    .Z(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06532_ (.I(_01352_),
    .Z(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06533_ (.I(_01353_),
    .Z(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06534_ (.I(_00654_),
    .ZN(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06535_ (.I(_01355_),
    .Z(_01356_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06536_ (.A1(_00700_),
    .A2(_00703_),
    .ZN(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06537_ (.I(_01357_),
    .Z(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06538_ (.I(_01358_),
    .Z(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06539_ (.I(_00640_),
    .Z(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06540_ (.A1(_01360_),
    .A2(_00647_),
    .ZN(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06541_ (.A1(_00694_),
    .A2(_00697_),
    .ZN(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06542_ (.I(_01362_),
    .Z(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06543_ (.I(_01363_),
    .Z(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06544_ (.I(_01364_),
    .Z(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06545_ (.A1(_00711_),
    .A2(_00712_),
    .ZN(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06546_ (.I(_00683_),
    .Z(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06547_ (.A1(net32),
    .A2(_01367_),
    .Z(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06548_ (.A1(net44),
    .A2(_00664_),
    .B(_01368_),
    .ZN(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06549_ (.A1(\as2650.insin[2] ),
    .A2(_00714_),
    .ZN(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06550_ (.A1(_00714_),
    .A2(_01369_),
    .B(_01370_),
    .ZN(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06551_ (.A1(_01366_),
    .A2(_01371_),
    .ZN(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06552_ (.I(_01372_),
    .Z(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06553_ (.I(_01373_),
    .Z(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06554_ (.I(_01374_),
    .Z(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06555_ (.I(_01375_),
    .Z(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06556_ (.I(_00708_),
    .Z(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06557_ (.A1(_00689_),
    .A2(_00693_),
    .ZN(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06558_ (.I(_01378_),
    .Z(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06559_ (.A1(_01377_),
    .A2(_01379_),
    .ZN(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06560_ (.A1(_01376_),
    .A2(_01380_),
    .ZN(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06561_ (.A1(_01365_),
    .A2(_01381_),
    .ZN(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06562_ (.A1(_01361_),
    .A2(_01382_),
    .ZN(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06563_ (.A1(_01359_),
    .A2(_01383_),
    .ZN(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06564_ (.I(_00643_),
    .Z(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06565_ (.A1(_01355_),
    .A2(_01385_),
    .A3(_00930_),
    .ZN(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06566_ (.I(_01386_),
    .Z(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06567_ (.A1(_00954_),
    .A2(_01387_),
    .ZN(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06568_ (.A1(_00679_),
    .A2(_00686_),
    .ZN(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06569_ (.A1(_01357_),
    .A2(_01389_),
    .ZN(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06570_ (.I(_01038_),
    .Z(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06571_ (.I(_01391_),
    .Z(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06572_ (.I(_01392_),
    .Z(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06573_ (.A1(_00713_),
    .A2(_00717_),
    .ZN(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06574_ (.I(_01394_),
    .Z(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06575_ (.I(_01395_),
    .Z(_01396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06576_ (.I(_01396_),
    .Z(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06577_ (.I(_01397_),
    .Z(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06578_ (.A1(_00698_),
    .A2(_01393_),
    .A3(_01398_),
    .ZN(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06579_ (.I(_01377_),
    .Z(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06580_ (.A1(_00675_),
    .A2(_00678_),
    .ZN(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06581_ (.A1(_00705_),
    .A2(_00706_),
    .ZN(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06582_ (.A1(_01401_),
    .A2(_01402_),
    .ZN(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06583_ (.A1(_01400_),
    .A2(_01403_),
    .ZN(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06584_ (.A1(_01399_),
    .A2(_01404_),
    .ZN(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06585_ (.I(_00713_),
    .Z(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06586_ (.A1(_00720_),
    .A2(_00721_),
    .ZN(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06587_ (.I(_01407_),
    .Z(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06588_ (.A1(_01400_),
    .A2(_01406_),
    .B(_01408_),
    .ZN(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06589_ (.A1(_01364_),
    .A2(_01390_),
    .A3(_01405_),
    .A4(_01409_),
    .ZN(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06590_ (.I(_01410_),
    .Z(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06591_ (.I(_01411_),
    .Z(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06592_ (.A1(_01224_),
    .A2(_01388_),
    .B(_01412_),
    .ZN(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06593_ (.A1(_01356_),
    .A2(_01384_),
    .B(_01413_),
    .ZN(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06594_ (.A1(_01245_),
    .A2(_01348_),
    .B(_01354_),
    .C(_01414_),
    .ZN(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06595_ (.I(_01415_),
    .ZN(net122));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06596_ (.I(_01367_),
    .Z(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06597_ (.I(_01416_),
    .Z(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06598_ (.I(_01417_),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06599_ (.A1(\as2650.ext_io_addr[7] ),
    .A2(\as2650.ext_io_addr[6] ),
    .ZN(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06600_ (.I(_01418_),
    .Z(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06601_ (.A1(\as2650.io_bus_we ),
    .A2(_01419_),
    .Z(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06602_ (.I(_01420_),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06603_ (.I(\as2650.ext_io_addr[6] ),
    .ZN(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06604_ (.A1(\as2650.ext_io_addr[7] ),
    .A2(_01421_),
    .ZN(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06605_ (.I(_01422_),
    .Z(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06606_ (.A1(\as2650.io_bus_we ),
    .A2(_01423_),
    .Z(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06607_ (.I(_01424_),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06608_ (.A1(\as2650.ext_io_addr[7] ),
    .A2(_01421_),
    .Z(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06609_ (.I(_01425_),
    .Z(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06610_ (.A1(\as2650.io_bus_we ),
    .A2(_01426_),
    .Z(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06611_ (.I(_01427_),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06612_ (.A1(\as2650.warmup[0] ),
    .A2(\as2650.warmup[1] ),
    .A3(net206),
    .ZN(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06613_ (.I(_01428_),
    .Z(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06614_ (.I(_01429_),
    .Z(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06615_ (.I(_01430_),
    .Z(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06616_ (.I(_01431_),
    .Z(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06617_ (.I(_01432_),
    .Z(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06618_ (.I(_01433_),
    .Z(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06619_ (.I(_01434_),
    .Z(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06620_ (.I(_01248_),
    .Z(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06621_ (.I(_01384_),
    .Z(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _06622_ (.A1(_01436_),
    .A2(_01318_),
    .A3(_01437_),
    .A4(net252),
    .Z(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06623_ (.A1(_01435_),
    .A2(_01438_),
    .ZN(net147));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06624_ (.A1(_01243_),
    .A2(_00956_),
    .ZN(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06625_ (.I(_01347_),
    .Z(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06626_ (.I(_01401_),
    .Z(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06627_ (.I(_01441_),
    .Z(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06628_ (.I(_01442_),
    .Z(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06629_ (.I(_01443_),
    .Z(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _06630_ (.A1(_01439_),
    .A2(_01440_),
    .B1(_01383_),
    .B2(_01444_),
    .ZN(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06631_ (.I(_01354_),
    .Z(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06632_ (.A1(_01446_),
    .A2(_01413_),
    .ZN(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06633_ (.A1(_01445_),
    .A2(_01447_),
    .ZN(net159));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06634_ (.I(_01431_),
    .Z(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06635_ (.I(_01448_),
    .Z(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06636_ (.I(_01449_),
    .Z(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06637_ (.A1(clknet_leaf_66_wb_clk_i),
    .A2(net204),
    .A3(_01450_),
    .Z(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06638_ (.I(_01451_),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06639_ (.A1(clknet_leaf_39_wb_clk_i),
    .A2(net205),
    .A3(_01450_),
    .Z(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06640_ (.I(_01452_),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06641_ (.A1(\web_behavior[1] ),
    .A2(clknet_leaf_159_wb_clk_i),
    .B(\web_behavior[0] ),
    .ZN(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06642_ (.A1(\web_behavior[1] ),
    .A2(clknet_leaf_159_wb_clk_i),
    .B(\web_behavior[0] ),
    .ZN(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06643__1 (.I(_01454_),
    .ZN(net292));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06644_ (.A1(_01453_),
    .A2(net292),
    .B(net252),
    .ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06645_ (.I(wb_debug_carry),
    .Z(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06646_ (.I(\as2650.debug_psl[0] ),
    .ZN(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06647_ (.I(_01457_),
    .Z(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06648_ (.I(\as2650.debug_psl[6] ),
    .Z(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06649_ (.I(_01459_),
    .Z(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06650_ (.I(_01402_),
    .Z(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06651_ (.I(_01461_),
    .Z(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06652_ (.A1(wb_debug_cc),
    .A2(_01245_),
    .ZN(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06653_ (.A1(wb_debug_cc),
    .A2(_01460_),
    .B1(_01462_),
    .B2(_01463_),
    .C(_01456_),
    .ZN(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06654_ (.A1(_01456_),
    .A2(_01458_),
    .B(_01464_),
    .ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06655_ (.I(\as2650.debug_psl[5] ),
    .ZN(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06656_ (.I(_01465_),
    .Z(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06657_ (.I(\as2650.debug_psl[7] ),
    .Z(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06658_ (.I(_01467_),
    .Z(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06659_ (.I(_01389_),
    .Z(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06660_ (.I(_01469_),
    .Z(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06661_ (.I(_01470_),
    .Z(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06662_ (.A1(wb_debug_cc),
    .A2(_01468_),
    .B1(_01471_),
    .B2(_01463_),
    .C(wb_debug_carry),
    .ZN(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06663_ (.A1(_01456_),
    .A2(_01466_),
    .B(_01472_),
    .ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06664_ (.I(_00583_),
    .Z(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06665_ (.I(_01473_),
    .Z(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06666_ (.I(_01474_),
    .Z(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06667_ (.I(_01475_),
    .Z(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06668_ (.I(_01476_),
    .Z(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06669_ (.I(_01477_),
    .Z(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06670_ (.I(_01478_),
    .Z(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06671_ (.I(_01479_),
    .Z(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06672_ (.I(_01478_),
    .Z(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06673_ (.A1(_01481_),
    .A2(\as2650.regs[6][0] ),
    .ZN(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06674_ (.A1(_01480_),
    .A2(_00869_),
    .B(_01482_),
    .ZN(net178));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06675_ (.A1(_01481_),
    .A2(\as2650.regs[6][1] ),
    .ZN(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06676_ (.A1(_01480_),
    .A2(_00854_),
    .B(_01483_),
    .ZN(net179));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06677_ (.I(_01478_),
    .Z(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06678_ (.A1(_01484_),
    .A2(\as2650.regs[6][2] ),
    .ZN(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06679_ (.A1(_01480_),
    .A2(_00897_),
    .B(_01485_),
    .ZN(net180));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06680_ (.A1(_01484_),
    .A2(\as2650.regs[6][3] ),
    .ZN(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06681_ (.A1(_01480_),
    .A2(_00884_),
    .B(_01486_),
    .ZN(net181));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06682_ (.A1(_01484_),
    .A2(\as2650.regs[6][4] ),
    .ZN(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06683_ (.A1(_01481_),
    .A2(_00837_),
    .B(_01487_),
    .ZN(net183));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06684_ (.A1(_01484_),
    .A2(\as2650.regs[6][5] ),
    .ZN(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06685_ (.A1(_01481_),
    .A2(_00818_),
    .B(_01488_),
    .ZN(net184));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06686_ (.I0(\as2650.regs[2][6] ),
    .I1(\as2650.regs[6][6] ),
    .S(_01479_),
    .Z(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06687_ (.I(_01489_),
    .Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06688_ (.I0(\as2650.regs[2][7] ),
    .I1(\as2650.regs[6][7] ),
    .S(_01479_),
    .Z(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06689_ (.I(_01490_),
    .Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06690_ (.I(_01473_),
    .Z(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06691_ (.A1(_01473_),
    .A2(\as2650.regs[7][0] ),
    .ZN(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06692_ (.A1(_01491_),
    .A2(_00999_),
    .B(_01492_),
    .ZN(net187));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06693_ (.A1(_01491_),
    .A2(\as2650.regs[7][1] ),
    .ZN(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06694_ (.A1(_01491_),
    .A2(_01017_),
    .B(_01493_),
    .ZN(net188));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06695_ (.A1(_01474_),
    .A2(\as2650.regs[7][2] ),
    .ZN(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06696_ (.A1(_01474_),
    .A2(_01040_),
    .B(_01494_),
    .ZN(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06697_ (.I(_01495_),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06698_ (.I0(\as2650.regs[3][3] ),
    .I1(\as2650.regs[7][3] ),
    .S(_01491_),
    .Z(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06699_ (.I(_01496_),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06700_ (.I(_00612_),
    .Z(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06701_ (.A1(_01497_),
    .A2(\as2650.regs[3][4] ),
    .ZN(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06702_ (.A1(_01497_),
    .A2(_00828_),
    .B(_01498_),
    .ZN(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06703_ (.I(_01499_),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06704_ (.A1(_00612_),
    .A2(\as2650.regs[3][5] ),
    .ZN(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06705_ (.A1(_00612_),
    .A2(_00810_),
    .B(_01500_),
    .ZN(net192));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06706_ (.I0(\as2650.regs[3][6] ),
    .I1(\as2650.regs[7][6] ),
    .S(_01475_),
    .Z(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06707_ (.I(_01501_),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06708_ (.I0(\as2650.regs[3][7] ),
    .I1(\as2650.regs[7][7] ),
    .S(_01474_),
    .Z(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06709_ (.I(_01502_),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06710_ (.I(_01377_),
    .Z(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06711_ (.I(_01503_),
    .Z(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06712_ (.I(_01504_),
    .Z(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06713_ (.A1(_00788_),
    .A2(_00912_),
    .ZN(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06714_ (.I(_01506_),
    .Z(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _06715_ (.A1(_00694_),
    .A2(_00697_),
    .Z(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06716_ (.A1(_01379_),
    .A2(_01508_),
    .ZN(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06717_ (.A1(_01375_),
    .A2(_01509_),
    .ZN(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06718_ (.A1(_01441_),
    .A2(_01461_),
    .A3(_01510_),
    .ZN(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06719_ (.A1(_01505_),
    .A2(_01507_),
    .A3(_01511_),
    .Z(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06720_ (.I(_01512_),
    .Z(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06721_ (.I(_00714_),
    .Z(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06722_ (.A1(_01514_),
    .A2(_01345_),
    .ZN(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06723_ (.A1(_01513_),
    .A2(_01515_),
    .ZN(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06724_ (.A1(\as2650.chirp_ptr[0] ),
    .A2(_01516_),
    .Z(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06725_ (.A1(_01352_),
    .A2(_01517_),
    .ZN(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06726_ (.I(_01518_),
    .Z(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06727_ (.I(\as2650.chirp_ptr[1] ),
    .ZN(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06728_ (.I(_01515_),
    .Z(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06729_ (.A1(\as2650.chirp_ptr[0] ),
    .A2(_01513_),
    .A3(_01520_),
    .ZN(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06730_ (.A1(_01519_),
    .A2(_01521_),
    .ZN(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06731_ (.A1(\as2650.chirp_ptr[2] ),
    .A2(_01522_),
    .Z(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06732_ (.I(_01523_),
    .ZN(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06733_ (.A1(_01432_),
    .A2(_01523_),
    .ZN(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06734_ (.I(_01525_),
    .ZN(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06735_ (.I(_01526_),
    .Z(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06736_ (.I(_00373_),
    .ZN(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06737_ (.A1(_01519_),
    .A2(_01521_),
    .Z(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06738_ (.A1(_01432_),
    .A2(_01528_),
    .ZN(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06739_ (.A1(_01527_),
    .A2(_01529_),
    .ZN(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06740_ (.A1(_01517_),
    .A2(_01529_),
    .Z(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06741_ (.A1(_01530_),
    .A2(_01531_),
    .ZN(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06742_ (.A1(_00373_),
    .A2(_01524_),
    .B1(_00375_),
    .B2(_01532_),
    .ZN(_00000_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06743_ (.A1(_01527_),
    .A2(_01525_),
    .A3(_01529_),
    .ZN(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06744_ (.A1(_01531_),
    .A2(_01533_),
    .ZN(_00001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06745_ (.A1(_01526_),
    .A2(_01528_),
    .ZN(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06746_ (.A1(_00375_),
    .A2(_01532_),
    .B(_01534_),
    .ZN(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06747_ (.A1(_01525_),
    .A2(_01531_),
    .ZN(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06748_ (.A1(_01526_),
    .A2(_01530_),
    .ZN(_00116_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06749_ (.A1(_01535_),
    .A2(_00116_),
    .Z(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06750_ (.I(_01536_),
    .Z(_00003_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06751_ (.A1(_01533_),
    .A2(_01534_),
    .Z(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06752_ (.I(_01537_),
    .Z(_00004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06753_ (.I(_01317_),
    .Z(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06754_ (.I(_01538_),
    .Z(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06755_ (.I(_01248_),
    .Z(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06756_ (.I(_01540_),
    .Z(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06757_ (.A1(_00661_),
    .A2(_00727_),
    .B(_01164_),
    .ZN(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06758_ (.A1(_01005_),
    .A2(_01542_),
    .ZN(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06759_ (.I(_00795_),
    .Z(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06760_ (.I(_00661_),
    .ZN(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06761_ (.A1(_00709_),
    .A2(_00718_),
    .A3(_00726_),
    .Z(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06762_ (.A1(_01545_),
    .A2(_01546_),
    .B(_01119_),
    .ZN(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06763_ (.A1(_01544_),
    .A2(_01320_),
    .ZN(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06764_ (.A1(_01544_),
    .A2(_01254_),
    .B(_01547_),
    .C(_01548_),
    .ZN(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _06765_ (.A1(_01543_),
    .A2(_01549_),
    .Z(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06766_ (.A1(_01211_),
    .A2(_01249_),
    .ZN(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06767_ (.A1(_01541_),
    .A2(_01550_),
    .B(_01551_),
    .ZN(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06768_ (.A1(_01539_),
    .A2(_01552_),
    .ZN(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06769_ (.I(_01318_),
    .Z(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06770_ (.A1(_01269_),
    .A2(_01554_),
    .ZN(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06771_ (.A1(_01553_),
    .A2(_01555_),
    .ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06772_ (.I(_01048_),
    .Z(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06773_ (.I(_01556_),
    .Z(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06774_ (.I(_01557_),
    .Z(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06775_ (.I(_01437_),
    .Z(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06776_ (.I(_01317_),
    .Z(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06777_ (.I(_01547_),
    .Z(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06778_ (.A1(_01023_),
    .A2(_01561_),
    .ZN(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06779_ (.I(_01542_),
    .Z(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _06780_ (.I(_01329_),
    .ZN(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06781_ (.A1(_01038_),
    .A2(_01564_),
    .ZN(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06782_ (.A1(_01391_),
    .A2(_01256_),
    .B(_01563_),
    .C(_01565_),
    .ZN(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06783_ (.A1(_01562_),
    .A2(_01566_),
    .ZN(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06784_ (.I(_01567_),
    .Z(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06785_ (.I0(_01207_),
    .I1(_01568_),
    .S(_01247_),
    .Z(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06786_ (.A1(_01560_),
    .A2(_01569_),
    .ZN(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06787_ (.I(_01318_),
    .Z(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06788_ (.I(_01384_),
    .Z(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06789_ (.A1(_01279_),
    .A2(_01571_),
    .B(_01572_),
    .ZN(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06790_ (.A1(_01558_),
    .A2(_01559_),
    .B1(_01570_),
    .B2(_01573_),
    .ZN(net167));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06791_ (.I(_01049_),
    .Z(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06792_ (.I(_01574_),
    .Z(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06793_ (.I(_01575_),
    .Z(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06794_ (.I(_01317_),
    .Z(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06795_ (.I(_01045_),
    .Z(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06796_ (.I(_00987_),
    .Z(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06797_ (.A1(_00987_),
    .A2(_01053_),
    .A3(_01054_),
    .ZN(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06798_ (.A1(_01579_),
    .A2(_01052_),
    .B(_01580_),
    .C(_01544_),
    .ZN(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06799_ (.A1(_01038_),
    .A2(_01333_),
    .B(_01547_),
    .ZN(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06800_ (.A1(_01578_),
    .A2(_01547_),
    .B1(_01581_),
    .B2(_01582_),
    .ZN(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06801_ (.A1(_01197_),
    .A2(_01248_),
    .ZN(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06802_ (.A1(_01249_),
    .A2(_01583_),
    .B(_01584_),
    .ZN(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06803_ (.A1(_01265_),
    .A2(_01538_),
    .ZN(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06804_ (.A1(_01577_),
    .A2(_01585_),
    .B(_01586_),
    .C(_01437_),
    .ZN(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06805_ (.A1(_01576_),
    .A2(_01559_),
    .B(_01587_),
    .ZN(net168));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06806_ (.I(_00974_),
    .Z(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06807_ (.I(_01588_),
    .Z(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06808_ (.I(_01589_),
    .Z(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06809_ (.I(_01339_),
    .ZN(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06810_ (.I(_01591_),
    .Z(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06811_ (.A1(_01391_),
    .A2(_01592_),
    .ZN(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06812_ (.A1(_01391_),
    .A2(_01070_),
    .A3(_01075_),
    .B(_01593_),
    .ZN(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06813_ (.I0(_01588_),
    .I1(_01594_),
    .S(_01563_),
    .Z(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06814_ (.I(_01595_),
    .Z(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06815_ (.A1(_01201_),
    .A2(_01540_),
    .ZN(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06816_ (.A1(_01436_),
    .A2(_01596_),
    .B(_01597_),
    .ZN(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06817_ (.A1(_01560_),
    .A2(_01598_),
    .ZN(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06818_ (.A1(_01287_),
    .A2(_01571_),
    .B(_01572_),
    .ZN(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06819_ (.A1(_01590_),
    .A2(_01559_),
    .B1(_01599_),
    .B2(_01600_),
    .ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06820_ (.I(_01089_),
    .Z(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06821_ (.I(_01601_),
    .Z(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06822_ (.I(_01602_),
    .Z(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06823_ (.A1(_01579_),
    .A2(_01098_),
    .B(_01101_),
    .ZN(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06824_ (.I(_01544_),
    .Z(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06825_ (.I0(_00638_),
    .I1(_01604_),
    .S(_01605_),
    .Z(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06826_ (.A1(_01089_),
    .A2(_01561_),
    .ZN(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06827_ (.A1(_01561_),
    .A2(_01606_),
    .B(_01607_),
    .ZN(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06828_ (.I(_01608_),
    .Z(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06829_ (.A1(_01162_),
    .A2(_01540_),
    .ZN(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06830_ (.A1(_01436_),
    .A2(_01609_),
    .B(_01610_),
    .ZN(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06831_ (.A1(_01577_),
    .A2(_01611_),
    .ZN(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06832_ (.A1(_01295_),
    .A2(_01554_),
    .B(_01572_),
    .ZN(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06833_ (.A1(_01603_),
    .A2(_01559_),
    .B1(_01612_),
    .B2(_01613_),
    .ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06834_ (.A1(_00813_),
    .A2(_00817_),
    .ZN(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06835_ (.A1(_00822_),
    .A2(_00826_),
    .ZN(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06836_ (.A1(_01614_),
    .A2(_01615_),
    .ZN(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06837_ (.I(_01561_),
    .Z(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06838_ (.I(_01605_),
    .Z(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06839_ (.A1(_00984_),
    .A2(_01090_),
    .ZN(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06840_ (.I0(_01088_),
    .I1(_01619_),
    .S(_01579_),
    .Z(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06841_ (.A1(_01618_),
    .A2(_01620_),
    .ZN(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06842_ (.I(_00627_),
    .Z(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06843_ (.A1(_01622_),
    .A2(_01392_),
    .B(_01617_),
    .ZN(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06844_ (.A1(_01616_),
    .A2(_01617_),
    .B1(_01621_),
    .B2(_01623_),
    .ZN(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06845_ (.I(_01624_),
    .Z(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06846_ (.A1(_01184_),
    .A2(_01249_),
    .ZN(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06847_ (.A1(_01541_),
    .A2(_01625_),
    .B(_01626_),
    .ZN(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06848_ (.A1(_01539_),
    .A2(_01627_),
    .ZN(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06849_ (.A1(_01301_),
    .A2(_01538_),
    .Z(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06850_ (.A1(_01628_),
    .A2(_01629_),
    .ZN(net154));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06851_ (.I(_00981_),
    .Z(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06852_ (.I(_01247_),
    .Z(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06853_ (.A1(_01239_),
    .A2(_01631_),
    .ZN(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06854_ (.I(_00917_),
    .Z(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06855_ (.I(_01617_),
    .Z(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06856_ (.A1(_00623_),
    .A2(_01605_),
    .ZN(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _06857_ (.A1(_01605_),
    .A2(_00988_),
    .B(_01617_),
    .C(_01635_),
    .ZN(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06858_ (.A1(_01633_),
    .A2(_01634_),
    .B(_01636_),
    .ZN(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06859_ (.I(_01637_),
    .Z(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06860_ (.A1(_01436_),
    .A2(_01638_),
    .ZN(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06861_ (.A1(_01632_),
    .A2(_01639_),
    .B(_01577_),
    .ZN(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06862_ (.A1(_01308_),
    .A2(_01554_),
    .B(_01437_),
    .ZN(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06863_ (.A1(_01630_),
    .A2(_01572_),
    .B1(_01640_),
    .B2(_01641_),
    .ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06864_ (.A1(_00907_),
    .A2(_00923_),
    .Z(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06865_ (.A1(_01392_),
    .A2(_01642_),
    .Z(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06866_ (.I(_00614_),
    .Z(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06867_ (.A1(_01644_),
    .A2(_01392_),
    .B(_01634_),
    .ZN(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06868_ (.A1(_00781_),
    .A2(_01634_),
    .B1(_01643_),
    .B2(_01645_),
    .ZN(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06869_ (.I(_01646_),
    .Z(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06870_ (.A1(_01214_),
    .A2(_01234_),
    .B(_01540_),
    .ZN(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06871_ (.A1(_01541_),
    .A2(_01647_),
    .B(_01648_),
    .ZN(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06872_ (.A1(_01539_),
    .A2(_01649_),
    .ZN(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06873_ (.A1(_01313_),
    .A2(_01554_),
    .ZN(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06874_ (.A1(_01650_),
    .A2(_01651_),
    .ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _06875_ (.A1(_01186_),
    .A2(_01213_),
    .A3(_01241_),
    .A4(_01315_),
    .Z(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06876_ (.I(_01652_),
    .Z(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06877_ (.I(_01653_),
    .Z(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06878_ (.I(_01654_),
    .Z(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06879_ (.A1(_01655_),
    .A2(_01387_),
    .ZN(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06880_ (.I(_01406_),
    .Z(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06881_ (.A1(_01377_),
    .A2(_01371_),
    .ZN(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06882_ (.I(_01658_),
    .Z(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06883_ (.A1(_01657_),
    .A2(_01659_),
    .ZN(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06884_ (.A1(_00658_),
    .A2(_01660_),
    .ZN(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06885_ (.I(_01371_),
    .Z(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06886_ (.A1(_01657_),
    .A2(_01662_),
    .B(_00954_),
    .ZN(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06887_ (.A1(_01661_),
    .A2(_01663_),
    .ZN(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06888_ (.A1(_01664_),
    .A2(_01656_),
    .ZN(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06889_ (.I(net296),
    .Z(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06890_ (.I(_01666_),
    .Z(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06891_ (.A1(net28),
    .A2(_00664_),
    .B(_00670_),
    .ZN(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06892_ (.I(_01668_),
    .Z(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06893_ (.A1(_01653_),
    .A2(_01428_),
    .A3(_01386_),
    .ZN(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06894_ (.I(_01670_),
    .Z(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06895_ (.A1(\as2650.instruction_args_latch[15] ),
    .A2(_01670_),
    .ZN(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06896_ (.A1(_01669_),
    .A2(_01671_),
    .B(_01672_),
    .ZN(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06897_ (.A1(_01228_),
    .A2(_01673_),
    .ZN(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06898_ (.A1(_01657_),
    .A2(_01662_),
    .ZN(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06899_ (.A1(_01674_),
    .A2(_01675_),
    .ZN(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06900_ (.A1(_01408_),
    .A2(_01676_),
    .ZN(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06901_ (.A1(_01667_),
    .A2(_01677_),
    .ZN(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06902_ (.I(_01656_),
    .Z(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06903_ (.I(_01679_),
    .Z(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06904_ (.I(_01680_),
    .Z(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06905_ (.A1(_00954_),
    .A2(_01514_),
    .A3(_01681_),
    .ZN(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06906_ (.I(_01353_),
    .Z(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06907_ (.I(_01683_),
    .Z(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06908_ (.I(_01684_),
    .Z(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06909_ (.A1(_01678_),
    .A2(_01682_),
    .B(_01685_),
    .ZN(_00005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06910_ (.I(net50),
    .Z(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06911_ (.I(net54),
    .Z(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06912_ (.I(net53),
    .Z(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06913_ (.A1(_01686_),
    .A2(_01687_),
    .A3(_01688_),
    .ZN(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06914_ (.A1(net88),
    .A2(net55),
    .ZN(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06915_ (.A1(wb_feedback_delay),
    .A2(_01690_),
    .ZN(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06916_ (.A1(net89),
    .A2(_01691_),
    .ZN(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _06917_ (.I(net51),
    .ZN(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06918_ (.A1(_01693_),
    .A2(net52),
    .ZN(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06919_ (.A1(_01692_),
    .A2(_01694_),
    .ZN(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06920_ (.A1(_01689_),
    .A2(_01695_),
    .ZN(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06921_ (.I(_01696_),
    .Z(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06922_ (.I(_01697_),
    .Z(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06923_ (.I0(net56),
    .I1(net106),
    .S(_01698_),
    .Z(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06924_ (.I(_01699_),
    .Z(_00006_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06925_ (.I0(net67),
    .I1(net113),
    .S(_01698_),
    .Z(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06926_ (.I(_01700_),
    .Z(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06927_ (.I0(net78),
    .I1(net114),
    .S(_01698_),
    .Z(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06928_ (.I(_01701_),
    .Z(_00008_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06929_ (.I0(net81),
    .I1(net115),
    .S(_01698_),
    .Z(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06930_ (.I(_01702_),
    .Z(_00009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06931_ (.I(_01697_),
    .Z(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06932_ (.I0(net82),
    .I1(net116),
    .S(_01703_),
    .Z(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06933_ (.I(_01704_),
    .Z(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06934_ (.I0(net83),
    .I1(net117),
    .S(_01703_),
    .Z(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06935_ (.I(_01705_),
    .Z(_00011_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06936_ (.I0(net84),
    .I1(net118),
    .S(_01703_),
    .Z(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06937_ (.I(_01706_),
    .Z(_00012_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06938_ (.I0(net85),
    .I1(net119),
    .S(_01703_),
    .Z(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06939_ (.I(_01707_),
    .Z(_00013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06940_ (.I(_01697_),
    .Z(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06941_ (.I0(net86),
    .I1(net120),
    .S(_01708_),
    .Z(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06942_ (.I(_01709_),
    .Z(_00014_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06943_ (.I0(net87),
    .I1(net121),
    .S(_01708_),
    .Z(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06944_ (.I(_01710_),
    .Z(_00015_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06945_ (.I0(net57),
    .I1(net107),
    .S(_01708_),
    .Z(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06946_ (.I(_01711_),
    .Z(_00016_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06947_ (.I0(net58),
    .I1(net108),
    .S(_01708_),
    .Z(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06948_ (.I(_01712_),
    .Z(_00017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06949_ (.I(_01697_),
    .Z(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06950_ (.I0(net59),
    .I1(net109),
    .S(_01713_),
    .Z(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06951_ (.I(_01714_),
    .Z(_00018_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06952_ (.I0(net60),
    .I1(net110),
    .S(_01713_),
    .Z(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06953_ (.I(_01715_),
    .Z(_00019_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06954_ (.I0(net61),
    .I1(net111),
    .S(_01713_),
    .Z(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06955_ (.I(_01716_),
    .Z(_00020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06956_ (.I0(net62),
    .I1(net112),
    .S(_01713_),
    .Z(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06957_ (.I(_01717_),
    .Z(_00021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06958_ (.I(_01696_),
    .Z(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06959_ (.I(_01718_),
    .Z(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06960_ (.I0(net63),
    .I1(net90),
    .S(_01719_),
    .Z(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06961_ (.I(_01720_),
    .Z(_00022_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06962_ (.I0(net64),
    .I1(net97),
    .S(_01719_),
    .Z(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06963_ (.I(_01721_),
    .Z(_00023_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06964_ (.I0(net65),
    .I1(net98),
    .S(_01719_),
    .Z(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06965_ (.I(_01722_),
    .Z(_00024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06966_ (.I0(net66),
    .I1(net99),
    .S(_01719_),
    .Z(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06967_ (.I(_01723_),
    .Z(_00025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06968_ (.I(_01718_),
    .Z(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06969_ (.I0(net68),
    .I1(net100),
    .S(_01724_),
    .Z(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06970_ (.I(_01725_),
    .Z(_00026_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06971_ (.I0(net69),
    .I1(net101),
    .S(_01724_),
    .Z(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06972_ (.I(_01726_),
    .Z(_00027_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06973_ (.I0(net70),
    .I1(net102),
    .S(_01724_),
    .Z(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06974_ (.I(_01727_),
    .Z(_00028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06975_ (.I0(net71),
    .I1(net103),
    .S(_01724_),
    .Z(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06976_ (.I(_01728_),
    .Z(_00029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06977_ (.I(_01718_),
    .Z(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06978_ (.I0(net72),
    .I1(net104),
    .S(_01729_),
    .Z(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06979_ (.I(_01730_),
    .Z(_00030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06980_ (.I0(net73),
    .I1(net105),
    .S(_01729_),
    .Z(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06981_ (.I(_01731_),
    .Z(_00031_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06982_ (.I0(net74),
    .I1(net91),
    .S(_01729_),
    .Z(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06983_ (.I(_01732_),
    .Z(_00032_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06984_ (.I0(net75),
    .I1(net92),
    .S(_01729_),
    .Z(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06985_ (.I(_01733_),
    .Z(_00033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06986_ (.I(_01718_),
    .Z(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06987_ (.I0(net76),
    .I1(net93),
    .S(_01734_),
    .Z(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06988_ (.I(_01735_),
    .Z(_00034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06989_ (.I0(net77),
    .I1(net94),
    .S(_01734_),
    .Z(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06990_ (.I(_01736_),
    .Z(_00035_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06991_ (.I0(net79),
    .I1(net95),
    .S(_01734_),
    .Z(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06992_ (.I(_01737_),
    .Z(_00036_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06993_ (.I0(net80),
    .I1(net96),
    .S(_01734_),
    .Z(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06994_ (.I(_01738_),
    .Z(_00037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06995_ (.I(_01686_),
    .Z(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06996_ (.I(net54),
    .Z(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06997_ (.I(_01740_),
    .Z(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06998_ (.I(net51),
    .Z(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06999_ (.I(net52),
    .Z(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07000_ (.I(_01688_),
    .ZN(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07001_ (.A1(_01687_),
    .A2(_01692_),
    .ZN(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07002_ (.A1(_01742_),
    .A2(_01743_),
    .A3(_01744_),
    .A4(_01745_),
    .ZN(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07003_ (.A1(_01739_),
    .A2(_01741_),
    .A3(net372),
    .ZN(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07004_ (.I0(net142),
    .I1(net56),
    .S(_01747_),
    .Z(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07005_ (.I(_01748_),
    .Z(_00038_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07006_ (.I0(net143),
    .I1(net67),
    .S(_01747_),
    .Z(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07007_ (.I(_01749_),
    .Z(_00039_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07008_ (.I0(net144),
    .I1(net78),
    .S(_01747_),
    .Z(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07009_ (.I(_01750_),
    .Z(_00040_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07010_ (.I(_01686_),
    .ZN(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07011_ (.I(_01751_),
    .Z(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07012_ (.I(_01752_),
    .Z(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07013_ (.A1(_01753_),
    .A2(wb_feedback_delay),
    .Z(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07014_ (.I(_01754_),
    .Z(_00041_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07015_ (.A1(wb_feedback_delay),
    .A2(_01690_),
    .Z(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07016_ (.I(_01755_),
    .Z(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07017_ (.I(_01756_),
    .Z(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07018_ (.A1(net216),
    .A2(_01757_),
    .ZN(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07019_ (.I(_01740_),
    .Z(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07020_ (.I(_01759_),
    .Z(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07021_ (.I(net53),
    .Z(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07022_ (.I(_01761_),
    .Z(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07023_ (.A1(_01693_),
    .A2(net106),
    .ZN(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07024_ (.A1(_01743_),
    .A2(_01744_),
    .ZN(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07025_ (.A1(_01742_),
    .A2(net142),
    .B(_01764_),
    .ZN(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07026_ (.A1(_01762_),
    .A2(_01458_),
    .B1(_01763_),
    .B2(_01765_),
    .ZN(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07027_ (.I(_01741_),
    .Z(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07028_ (.I(\wb_counter[0] ),
    .ZN(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07029_ (.A1(_01767_),
    .A2(_01768_),
    .ZN(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07030_ (.I(_01691_),
    .Z(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07031_ (.A1(_01760_),
    .A2(_01766_),
    .B(_01769_),
    .C(_01770_),
    .ZN(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07032_ (.I(_01739_),
    .Z(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07033_ (.I(_01772_),
    .Z(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07034_ (.A1(_01758_),
    .A2(_01771_),
    .B(_01773_),
    .ZN(_00042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07035_ (.A1(net227),
    .A2(_01757_),
    .ZN(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _07036_ (.I(\as2650.debug_psl[1] ),
    .ZN(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07037_ (.A1(_01693_),
    .A2(net113),
    .ZN(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07038_ (.A1(_01742_),
    .A2(net143),
    .B(_01764_),
    .ZN(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07039_ (.A1(_01762_),
    .A2(_01775_),
    .B1(_01776_),
    .B2(_01777_),
    .ZN(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07040_ (.I(_01687_),
    .Z(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07041_ (.I(_01779_),
    .Z(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07042_ (.I(\wb_counter[1] ),
    .ZN(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07043_ (.A1(_01780_),
    .A2(_01781_),
    .ZN(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07044_ (.A1(_01760_),
    .A2(_01778_),
    .B(_01782_),
    .C(_01770_),
    .ZN(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07045_ (.A1(_01774_),
    .A2(_01783_),
    .B(_01773_),
    .ZN(_00043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07046_ (.A1(net238),
    .A2(_01757_),
    .ZN(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _07047_ (.I(\as2650.debug_psl[2] ),
    .ZN(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07048_ (.A1(_01693_),
    .A2(net114),
    .ZN(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07049_ (.A1(_01742_),
    .A2(net144),
    .B(_01764_),
    .ZN(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07050_ (.A1(_01762_),
    .A2(_01785_),
    .B1(_01786_),
    .B2(_01787_),
    .ZN(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07051_ (.I(\wb_counter[2] ),
    .ZN(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07052_ (.A1(_01780_),
    .A2(_01789_),
    .ZN(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07053_ (.A1(_01760_),
    .A2(_01788_),
    .B(_01790_),
    .C(_01770_),
    .ZN(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07054_ (.A1(_01784_),
    .A2(_01791_),
    .B(_01773_),
    .ZN(_00044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07055_ (.I(_01686_),
    .Z(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07056_ (.I(_01792_),
    .Z(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07057_ (.I(_01755_),
    .Z(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07058_ (.I(_01794_),
    .Z(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07059_ (.I(\wb_counter[3] ),
    .ZN(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07060_ (.I(net357),
    .Z(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07061_ (.I(_01797_),
    .Z(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07062_ (.A1(net51),
    .A2(_01743_),
    .B(_01688_),
    .ZN(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07063_ (.I(_01799_),
    .Z(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07064_ (.A1(net115),
    .A2(_01798_),
    .B(_01800_),
    .ZN(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07065_ (.I(\as2650.debug_psl[3] ),
    .Z(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07066_ (.I(_01802_),
    .Z(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07067_ (.I(_01803_),
    .Z(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07068_ (.I(_01740_),
    .Z(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07069_ (.A1(_01762_),
    .A2(_01804_),
    .B(_01805_),
    .ZN(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07070_ (.I(_01755_),
    .Z(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07071_ (.I(_01807_),
    .Z(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07072_ (.A1(_01780_),
    .A2(_01796_),
    .B1(_01801_),
    .B2(_01806_),
    .C(_01808_),
    .ZN(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07073_ (.A1(net241),
    .A2(_01795_),
    .B(_01809_),
    .ZN(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07074_ (.A1(_01793_),
    .A2(_01810_),
    .ZN(_00045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07075_ (.I(\wb_counter[4] ),
    .ZN(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07076_ (.A1(net116),
    .A2(_01798_),
    .B(_01800_),
    .ZN(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07077_ (.I(_01475_),
    .Z(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07078_ (.I(_01813_),
    .Z(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07079_ (.I(_01688_),
    .Z(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07080_ (.I(_01779_),
    .Z(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07081_ (.A1(_01814_),
    .A2(_01815_),
    .B(_01816_),
    .ZN(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07082_ (.A1(_01780_),
    .A2(_01811_),
    .B1(_01812_),
    .B2(_01817_),
    .C(_01808_),
    .ZN(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07083_ (.A1(net242),
    .A2(_01795_),
    .B(_01818_),
    .ZN(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07084_ (.A1(_01793_),
    .A2(_01819_),
    .ZN(_00046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07085_ (.I(_01739_),
    .Z(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07086_ (.I(_01820_),
    .Z(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07087_ (.I(_01741_),
    .Z(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07088_ (.I(\wb_counter[5] ),
    .ZN(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07089_ (.A1(net117),
    .A2(_01798_),
    .B(_01800_),
    .ZN(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07090_ (.I(_01761_),
    .Z(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07091_ (.I(\as2650.debug_psl[5] ),
    .Z(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07092_ (.I(_01826_),
    .Z(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07093_ (.A1(_01825_),
    .A2(_01827_),
    .B(_01816_),
    .ZN(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07094_ (.A1(_01822_),
    .A2(_01823_),
    .B1(_01824_),
    .B2(_01828_),
    .C(_01808_),
    .ZN(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07095_ (.A1(net243),
    .A2(_01795_),
    .B(_01829_),
    .ZN(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07096_ (.A1(_01821_),
    .A2(_01830_),
    .ZN(_00047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07097_ (.I(\wb_counter[6] ),
    .ZN(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07098_ (.A1(net118),
    .A2(_01798_),
    .B(_01800_),
    .ZN(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07099_ (.A1(_01460_),
    .A2(_01815_),
    .B(_01816_),
    .ZN(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07100_ (.A1(_01822_),
    .A2(_01831_),
    .B1(_01832_),
    .B2(_01833_),
    .C(_01808_),
    .ZN(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07101_ (.A1(net244),
    .A2(_01795_),
    .B(_01834_),
    .ZN(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07102_ (.A1(_01821_),
    .A2(_01835_),
    .ZN(_00048_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07103_ (.I(_01794_),
    .Z(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07104_ (.I(\wb_counter[7] ),
    .ZN(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07105_ (.I(_01797_),
    .Z(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07106_ (.I(_01799_),
    .Z(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07107_ (.A1(net119),
    .A2(_01838_),
    .B(_01839_),
    .ZN(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07108_ (.A1(_01468_),
    .A2(_01815_),
    .B(_01816_),
    .ZN(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07109_ (.I(_01807_),
    .Z(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07110_ (.A1(_01822_),
    .A2(_01837_),
    .B1(_01840_),
    .B2(_01841_),
    .C(_01842_),
    .ZN(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07111_ (.A1(net245),
    .A2(_01836_),
    .B(_01843_),
    .ZN(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07112_ (.A1(_01821_),
    .A2(_01844_),
    .ZN(_00049_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07113_ (.I(\wb_counter[8] ),
    .ZN(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07114_ (.A1(net120),
    .A2(_01838_),
    .B(_01839_),
    .ZN(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07115_ (.I(\as2650.debug_psu[0] ),
    .Z(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07116_ (.I(_01847_),
    .Z(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07117_ (.I(_01848_),
    .Z(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07118_ (.I(_01779_),
    .Z(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07119_ (.A1(_01825_),
    .A2(_01849_),
    .B(_01850_),
    .ZN(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07120_ (.A1(_01822_),
    .A2(_01845_),
    .B1(_01846_),
    .B2(_01851_),
    .C(_01842_),
    .ZN(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07121_ (.A1(net246),
    .A2(_01836_),
    .B(_01852_),
    .ZN(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07122_ (.A1(_01821_),
    .A2(_01853_),
    .ZN(_00050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07123_ (.I(_01772_),
    .Z(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07124_ (.I(_01741_),
    .Z(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07125_ (.I(\wb_counter[9] ),
    .ZN(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07126_ (.A1(net121),
    .A2(_01838_),
    .B(_01839_),
    .ZN(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07127_ (.I(\as2650.debug_psu[1] ),
    .Z(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07128_ (.I(_01858_),
    .Z(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07129_ (.I(_01859_),
    .Z(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07130_ (.A1(_01825_),
    .A2(_01860_),
    .B(_01850_),
    .ZN(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07131_ (.A1(_01855_),
    .A2(_01856_),
    .B1(_01857_),
    .B2(_01861_),
    .C(_01842_),
    .ZN(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07132_ (.A1(net247),
    .A2(_01836_),
    .B(_01862_),
    .ZN(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07133_ (.A1(_01854_),
    .A2(_01863_),
    .ZN(_00051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07134_ (.I(\wb_counter[10] ),
    .ZN(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07135_ (.A1(net107),
    .A2(_01838_),
    .B(_01839_),
    .ZN(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07136_ (.I(\as2650.debug_psu[2] ),
    .Z(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07137_ (.I(_01866_),
    .Z(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07138_ (.I(_01867_),
    .Z(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07139_ (.I(_01868_),
    .Z(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07140_ (.A1(_01825_),
    .A2(_01869_),
    .B(_01850_),
    .ZN(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07141_ (.A1(_01855_),
    .A2(_01864_),
    .B1(_01865_),
    .B2(_01870_),
    .C(_01842_),
    .ZN(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07142_ (.A1(net217),
    .A2(_01836_),
    .B(_01871_),
    .ZN(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07143_ (.A1(_01854_),
    .A2(_01872_),
    .ZN(_00052_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07144_ (.I(_01794_),
    .Z(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07145_ (.I(\wb_counter[11] ),
    .ZN(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07146_ (.I(_01797_),
    .Z(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07147_ (.I(_01799_),
    .Z(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07148_ (.A1(net108),
    .A2(_01875_),
    .B(_01876_),
    .ZN(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07149_ (.I(_01761_),
    .Z(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07150_ (.I(\as2650.debug_psu[3] ),
    .Z(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07151_ (.I(_01879_),
    .Z(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07152_ (.I(_01880_),
    .Z(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07153_ (.A1(_01878_),
    .A2(_01881_),
    .B(_01850_),
    .ZN(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07154_ (.I(_01755_),
    .Z(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07155_ (.A1(_01855_),
    .A2(_01874_),
    .B1(_01877_),
    .B2(_01882_),
    .C(_01883_),
    .ZN(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07156_ (.A1(net218),
    .A2(_01873_),
    .B(_01884_),
    .ZN(_01885_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07157_ (.A1(_01854_),
    .A2(_01885_),
    .ZN(_00053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07158_ (.I(\wb_counter[12] ),
    .ZN(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07159_ (.A1(net109),
    .A2(_01875_),
    .B(_01876_),
    .ZN(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07160_ (.I(\as2650.debug_psu[4] ),
    .Z(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07161_ (.I(_01740_),
    .Z(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07162_ (.A1(_01878_),
    .A2(_01888_),
    .B(_01889_),
    .ZN(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07163_ (.A1(_01855_),
    .A2(_01886_),
    .B1(_01887_),
    .B2(_01890_),
    .C(_01883_),
    .ZN(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07164_ (.A1(net219),
    .A2(_01873_),
    .B(_01891_),
    .ZN(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07165_ (.A1(_01854_),
    .A2(_01892_),
    .ZN(_00054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07166_ (.I(_01772_),
    .Z(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07167_ (.I(\wb_counter[13] ),
    .ZN(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07168_ (.A1(net110),
    .A2(_01875_),
    .B(_01876_),
    .ZN(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07169_ (.I(\as2650.debug_psu[5] ),
    .Z(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07170_ (.I(_01896_),
    .Z(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07171_ (.A1(_01878_),
    .A2(_01897_),
    .B(_01889_),
    .ZN(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07172_ (.A1(_01805_),
    .A2(_01894_),
    .B1(_01895_),
    .B2(_01898_),
    .C(_01883_),
    .ZN(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07173_ (.A1(net220),
    .A2(_01873_),
    .B(_01899_),
    .ZN(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07174_ (.A1(_01893_),
    .A2(_01900_),
    .ZN(_00055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07175_ (.I(\wb_counter[14] ),
    .ZN(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07176_ (.A1(net111),
    .A2(_01875_),
    .B(_01876_),
    .ZN(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07177_ (.I(net253),
    .Z(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07178_ (.A1(_01878_),
    .A2(_01903_),
    .B(_01889_),
    .ZN(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07179_ (.A1(_01805_),
    .A2(_01901_),
    .B1(_01902_),
    .B2(_01904_),
    .C(_01883_),
    .ZN(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07180_ (.A1(net221),
    .A2(_01873_),
    .B(_01905_),
    .ZN(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07181_ (.A1(_01893_),
    .A2(_01906_),
    .ZN(_00056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07182_ (.I(\wb_counter[15] ),
    .ZN(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07183_ (.I(net357),
    .Z(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07184_ (.A1(net112),
    .A2(_01908_),
    .B(_01799_),
    .ZN(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07185_ (.I(\as2650.debug_psu[7] ),
    .Z(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07186_ (.A1(_01815_),
    .A2(_01910_),
    .B(_01889_),
    .ZN(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07187_ (.A1(_01805_),
    .A2(_01907_),
    .B1(_01909_),
    .B2(_01911_),
    .C(_01794_),
    .ZN(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07188_ (.A1(net222),
    .A2(_01757_),
    .B(_01912_),
    .ZN(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07189_ (.A1(_01893_),
    .A2(_01913_),
    .ZN(_00057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07190_ (.I(net223),
    .ZN(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07191_ (.I(_01807_),
    .Z(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07192_ (.I(_01915_),
    .Z(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07193_ (.I(_01908_),
    .Z(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07194_ (.A1(net51),
    .A2(_01743_),
    .ZN(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07195_ (.A1(net346),
    .A2(net53),
    .ZN(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07196_ (.A1(_01918_),
    .A2(_01919_),
    .Z(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07197_ (.I(_01920_),
    .Z(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07198_ (.I(_01921_),
    .Z(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07199_ (.A1(net90),
    .A2(_01917_),
    .B(_01922_),
    .ZN(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07200_ (.I(_01756_),
    .Z(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07201_ (.A1(_01760_),
    .A2(\wb_counter[16] ),
    .B(_01924_),
    .ZN(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07202_ (.I(_01739_),
    .Z(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07203_ (.A1(_01914_),
    .A2(_01916_),
    .B1(_01923_),
    .B2(_01925_),
    .C(_01926_),
    .ZN(_00058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07204_ (.I(net224),
    .ZN(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07205_ (.A1(net97),
    .A2(_01917_),
    .B(_01922_),
    .ZN(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07206_ (.I(_01759_),
    .Z(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07207_ (.A1(_01929_),
    .A2(\wb_counter[17] ),
    .B(_01924_),
    .ZN(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07208_ (.I(_01792_),
    .Z(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07209_ (.A1(_01927_),
    .A2(_01916_),
    .B1(_01928_),
    .B2(_01930_),
    .C(_01931_),
    .ZN(_00059_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07210_ (.I(net225),
    .ZN(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07211_ (.A1(net98),
    .A2(_01917_),
    .B(_01922_),
    .ZN(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07212_ (.A1(_01929_),
    .A2(\wb_counter[18] ),
    .B(_01924_),
    .ZN(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07213_ (.A1(_01932_),
    .A2(_01916_),
    .B1(_01933_),
    .B2(_01934_),
    .C(_01931_),
    .ZN(_00060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07214_ (.I(net226),
    .ZN(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07215_ (.I(_01919_),
    .Z(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07216_ (.A1(net99),
    .A2(_01917_),
    .B(_01936_),
    .ZN(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07217_ (.A1(_01929_),
    .A2(\wb_counter[19] ),
    .B(_01924_),
    .ZN(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07218_ (.A1(_01935_),
    .A2(_01916_),
    .B1(_01937_),
    .B2(_01938_),
    .C(_01931_),
    .ZN(_00061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07219_ (.I(net228),
    .ZN(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07220_ (.I(_01915_),
    .Z(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07221_ (.I(_01908_),
    .Z(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07222_ (.A1(net100),
    .A2(_01941_),
    .B(_01922_),
    .ZN(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07223_ (.I(_01756_),
    .Z(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07224_ (.A1(_01929_),
    .A2(\wb_counter[20] ),
    .B(_01943_),
    .ZN(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07225_ (.A1(_01939_),
    .A2(_01940_),
    .B1(_01942_),
    .B2(_01944_),
    .C(_01931_),
    .ZN(_00062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07226_ (.I(net229),
    .ZN(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07227_ (.I(_01920_),
    .Z(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07228_ (.A1(net101),
    .A2(_01941_),
    .B(_01946_),
    .ZN(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07229_ (.I(_01759_),
    .Z(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07230_ (.A1(_01948_),
    .A2(\wb_counter[21] ),
    .B(_01943_),
    .ZN(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07231_ (.I(_01792_),
    .Z(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07232_ (.A1(_01945_),
    .A2(_01940_),
    .B1(_01947_),
    .B2(_01949_),
    .C(_01950_),
    .ZN(_00063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07233_ (.I(net230),
    .ZN(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07234_ (.A1(net102),
    .A2(_01941_),
    .B(_01946_),
    .ZN(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07235_ (.A1(_01948_),
    .A2(\wb_counter[22] ),
    .B(_01943_),
    .ZN(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07236_ (.A1(_01951_),
    .A2(_01940_),
    .B1(_01952_),
    .B2(_01953_),
    .C(_01950_),
    .ZN(_00064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07237_ (.I(net231),
    .ZN(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07238_ (.A1(net103),
    .A2(_01941_),
    .B(_01946_),
    .ZN(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07239_ (.A1(_01948_),
    .A2(\wb_counter[23] ),
    .B(_01943_),
    .ZN(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07240_ (.A1(_01954_),
    .A2(_01940_),
    .B1(_01955_),
    .B2(_01956_),
    .C(_01950_),
    .ZN(_00065_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07241_ (.I(net232),
    .ZN(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07242_ (.I(_01915_),
    .Z(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07243_ (.I(_01908_),
    .Z(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07244_ (.A1(net104),
    .A2(_01959_),
    .B(_01936_),
    .ZN(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07245_ (.I(_01756_),
    .Z(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07246_ (.A1(_01948_),
    .A2(\wb_counter[24] ),
    .B(_01961_),
    .ZN(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07247_ (.A1(_01957_),
    .A2(_01958_),
    .B1(_01960_),
    .B2(_01962_),
    .C(_01950_),
    .ZN(_00066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07248_ (.I(net233),
    .ZN(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07249_ (.A1(net105),
    .A2(_01959_),
    .B(_01946_),
    .ZN(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07250_ (.I(_01759_),
    .Z(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07251_ (.A1(_01965_),
    .A2(\wb_counter[25] ),
    .B(_01961_),
    .ZN(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07252_ (.I(_01792_),
    .Z(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07253_ (.A1(_01963_),
    .A2(_01958_),
    .B1(_01964_),
    .B2(_01966_),
    .C(_01967_),
    .ZN(_00067_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07254_ (.I(net234),
    .ZN(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07255_ (.A1(net91),
    .A2(_01959_),
    .B(_01921_),
    .ZN(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07256_ (.A1(_01965_),
    .A2(\wb_counter[26] ),
    .B(_01961_),
    .ZN(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07257_ (.A1(_01968_),
    .A2(_01958_),
    .B1(_01969_),
    .B2(_01970_),
    .C(_01967_),
    .ZN(_00068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07258_ (.I(net235),
    .ZN(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07259_ (.A1(net92),
    .A2(_01959_),
    .B(_01921_),
    .ZN(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07260_ (.A1(_01965_),
    .A2(\wb_counter[27] ),
    .B(_01961_),
    .ZN(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07261_ (.A1(_01971_),
    .A2(_01958_),
    .B1(_01972_),
    .B2(_01973_),
    .C(_01967_),
    .ZN(_00069_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07262_ (.I(net236),
    .ZN(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07263_ (.I(_01915_),
    .Z(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07264_ (.I(_01797_),
    .Z(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07265_ (.A1(net93),
    .A2(_01976_),
    .B(_01936_),
    .ZN(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07266_ (.I(_01807_),
    .Z(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07267_ (.A1(_01965_),
    .A2(\wb_counter[28] ),
    .B(_01978_),
    .ZN(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07268_ (.A1(_01974_),
    .A2(_01975_),
    .B1(_01977_),
    .B2(_01979_),
    .C(_01967_),
    .ZN(_00070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07269_ (.I(net237),
    .ZN(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07270_ (.A1(net94),
    .A2(_01976_),
    .B(_01936_),
    .ZN(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07271_ (.A1(_01767_),
    .A2(\wb_counter[29] ),
    .B(_01978_),
    .ZN(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07272_ (.A1(_01980_),
    .A2(_01975_),
    .B1(_01981_),
    .B2(_01982_),
    .C(_01820_),
    .ZN(_00071_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07273_ (.I(net239),
    .ZN(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07274_ (.A1(net95),
    .A2(_01976_),
    .B(_01921_),
    .ZN(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07275_ (.A1(_01767_),
    .A2(\wb_counter[30] ),
    .B(_01978_),
    .ZN(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07276_ (.A1(_01983_),
    .A2(_01975_),
    .B1(_01984_),
    .B2(_01985_),
    .C(_01820_),
    .ZN(_00072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07277_ (.I(net240),
    .ZN(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _07278_ (.A1(net96),
    .A2(_01976_),
    .B1(_01918_),
    .B2(_00684_),
    .C(_01919_),
    .ZN(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07279_ (.A1(_01767_),
    .A2(\wb_counter[31] ),
    .B(_01978_),
    .ZN(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07280_ (.A1(_01986_),
    .A2(_01975_),
    .B1(net392),
    .B2(_01988_),
    .C(_01820_),
    .ZN(_00073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07281_ (.A1(_01893_),
    .A2(net378),
    .ZN(_00074_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07282_ (.A1(_01779_),
    .A2(_01744_),
    .A3(_01692_),
    .ZN(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07283_ (.I(_01989_),
    .Z(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07284_ (.A1(net334),
    .A2(_01990_),
    .ZN(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07285_ (.A1(_01761_),
    .A2(_01745_),
    .ZN(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07286_ (.I(_01992_),
    .Z(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07287_ (.A1(wb_debug_cc),
    .A2(_01993_),
    .ZN(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07288_ (.A1(net335),
    .A2(_01994_),
    .B(_01773_),
    .ZN(_00075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07289_ (.A1(net67),
    .A2(_01990_),
    .ZN(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07290_ (.A1(_01456_),
    .A2(_01993_),
    .ZN(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07291_ (.I(_01772_),
    .Z(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07292_ (.A1(net348),
    .A2(_01996_),
    .B(_01997_),
    .ZN(_00076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07293_ (.A1(net312),
    .A2(_01990_),
    .ZN(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07294_ (.A1(\web_behavior[0] ),
    .A2(_01993_),
    .ZN(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07295_ (.A1(net313),
    .A2(_01999_),
    .B(_01997_),
    .ZN(_00077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07296_ (.A1(net304),
    .A2(_01990_),
    .ZN(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07297_ (.I(_01992_),
    .Z(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07298_ (.A1(\web_behavior[1] ),
    .A2(_02001_),
    .ZN(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07299_ (.A1(net305),
    .A2(_02002_),
    .B(_01997_),
    .ZN(_00078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07300_ (.A1(net82),
    .A2(_01989_),
    .ZN(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07301_ (.A1(wb_reset_override_en),
    .A2(_02001_),
    .ZN(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07302_ (.A1(net316),
    .A2(_02004_),
    .B(_01997_),
    .ZN(_00079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07303_ (.A1(net83),
    .A2(_01989_),
    .ZN(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07304_ (.A1(wb_reset_override),
    .A2(_02001_),
    .ZN(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07305_ (.A1(net323),
    .A2(_02006_),
    .B(_01793_),
    .ZN(_00080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07306_ (.A1(net84),
    .A2(_01992_),
    .B(_01753_),
    .ZN(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07307_ (.A1(net148),
    .A2(_01993_),
    .B(_02007_),
    .ZN(_00081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07308_ (.A1(net85),
    .A2(_01989_),
    .ZN(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07309_ (.A1(net165),
    .A2(_02001_),
    .ZN(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07310_ (.A1(net319),
    .A2(_02009_),
    .B(_01793_),
    .ZN(_00082_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _07311_ (.I(_00684_),
    .ZN(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07312_ (.A1(net80),
    .A2(net372),
    .B(_01753_),
    .ZN(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07313_ (.A1(_02010_),
    .A2(net372),
    .B(_02011_),
    .ZN(_00083_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07314_ (.A1(net89),
    .A2(_01687_),
    .A3(_01770_),
    .ZN(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07315_ (.I(_02012_),
    .Z(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07316_ (.I(_02013_),
    .Z(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07317_ (.A1(net56),
    .A2(_02013_),
    .ZN(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07318_ (.A1(\wb_counter[0] ),
    .A2(_02014_),
    .B(_02015_),
    .C(_01926_),
    .ZN(_00084_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07319_ (.A1(_01768_),
    .A2(\wb_counter[1] ),
    .Z(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07320_ (.A1(net67),
    .A2(_02013_),
    .ZN(_02017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07321_ (.A1(_02014_),
    .A2(_02016_),
    .B(_02017_),
    .C(_01926_),
    .ZN(_00085_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07322_ (.A1(\wb_counter[0] ),
    .A2(\wb_counter[1] ),
    .A3(\wb_counter[2] ),
    .ZN(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07323_ (.A1(_01768_),
    .A2(_01781_),
    .B(_01789_),
    .ZN(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07324_ (.A1(_02018_),
    .A2(_02019_),
    .ZN(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07325_ (.A1(net78),
    .A2(_02013_),
    .ZN(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07326_ (.A1(_02014_),
    .A2(_02020_),
    .B(_02021_),
    .C(_01926_),
    .ZN(_00086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07327_ (.I(_02012_),
    .Z(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07328_ (.I(_02022_),
    .Z(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07329_ (.I(_02023_),
    .Z(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07330_ (.A1(\wb_counter[3] ),
    .A2(_02018_),
    .Z(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07331_ (.I(_02012_),
    .Z(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07332_ (.I(_02026_),
    .Z(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07333_ (.A1(net304),
    .A2(_02027_),
    .B(_01753_),
    .ZN(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07334_ (.A1(_02024_),
    .A2(_02025_),
    .B(_02028_),
    .ZN(_00087_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07335_ (.A1(_01796_),
    .A2(_02018_),
    .ZN(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07336_ (.A1(_01811_),
    .A2(_02029_),
    .Z(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07337_ (.I(_01752_),
    .Z(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07338_ (.A1(net82),
    .A2(_02027_),
    .B(_02031_),
    .ZN(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07339_ (.A1(_02024_),
    .A2(_02030_),
    .B(_02032_),
    .ZN(_00088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07340_ (.A1(\wb_counter[4] ),
    .A2(_02029_),
    .ZN(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07341_ (.A1(_01823_),
    .A2(_02033_),
    .ZN(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07342_ (.A1(\wb_counter[4] ),
    .A2(\wb_counter[5] ),
    .A3(_02029_),
    .ZN(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07343_ (.A1(_02034_),
    .A2(_02035_),
    .ZN(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07344_ (.A1(net322),
    .A2(_02027_),
    .B(_02031_),
    .ZN(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07345_ (.A1(_02024_),
    .A2(_02036_),
    .B(_02037_),
    .ZN(_00089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07346_ (.A1(_01831_),
    .A2(_02035_),
    .ZN(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07347_ (.A1(_01831_),
    .A2(_02035_),
    .Z(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07348_ (.A1(_02038_),
    .A2(_02039_),
    .ZN(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07349_ (.A1(net84),
    .A2(_02027_),
    .B(_02031_),
    .ZN(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07350_ (.A1(_02024_),
    .A2(_02040_),
    .B(_02041_),
    .ZN(_00090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07351_ (.I(_02023_),
    .Z(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07352_ (.A1(\wb_counter[7] ),
    .A2(_02039_),
    .Z(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07353_ (.I(_02026_),
    .Z(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07354_ (.A1(net85),
    .A2(_02044_),
    .B(_02031_),
    .ZN(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07355_ (.A1(_02042_),
    .A2(_02043_),
    .B(_02045_),
    .ZN(_00091_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07356_ (.A1(_01837_),
    .A2(_02039_),
    .ZN(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07357_ (.A1(_01845_),
    .A2(_02046_),
    .Z(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07358_ (.I(_01752_),
    .Z(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07359_ (.A1(net338),
    .A2(_02044_),
    .B(_02048_),
    .ZN(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07360_ (.A1(_02042_),
    .A2(_02047_),
    .B(net339),
    .ZN(_00092_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07361_ (.A1(_01837_),
    .A2(_01845_),
    .A3(_02039_),
    .ZN(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07362_ (.A1(_01856_),
    .A2(_02050_),
    .Z(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07363_ (.A1(net326),
    .A2(_02044_),
    .B(_02048_),
    .ZN(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07364_ (.A1(_02042_),
    .A2(_02051_),
    .B(net327),
    .ZN(_00093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07365_ (.A1(\wb_counter[9] ),
    .A2(_02050_),
    .ZN(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07366_ (.A1(\wb_counter[10] ),
    .A2(_02053_),
    .Z(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07367_ (.A1(net330),
    .A2(_02044_),
    .B(_02048_),
    .ZN(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07368_ (.A1(_02042_),
    .A2(_02054_),
    .B(net331),
    .ZN(_00094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07369_ (.I(_02023_),
    .Z(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07370_ (.A1(_01864_),
    .A2(_02053_),
    .ZN(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07371_ (.A1(_01874_),
    .A2(_02057_),
    .Z(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07372_ (.I(_02026_),
    .Z(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07373_ (.A1(net342),
    .A2(_02059_),
    .B(_02048_),
    .ZN(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07374_ (.A1(_02056_),
    .A2(_02058_),
    .B(net343),
    .ZN(_00095_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07375_ (.A1(\wb_counter[11] ),
    .A2(\wb_counter[12] ),
    .A3(_02057_),
    .ZN(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07376_ (.A1(\wb_counter[11] ),
    .A2(_02057_),
    .ZN(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07377_ (.A1(_01886_),
    .A2(_02062_),
    .ZN(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07378_ (.A1(_02061_),
    .A2(_02063_),
    .ZN(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07379_ (.I(_01752_),
    .Z(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07380_ (.A1(net308),
    .A2(_02059_),
    .B(_02065_),
    .ZN(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07381_ (.A1(_02056_),
    .A2(_02064_),
    .B(net309),
    .ZN(_00096_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07382_ (.A1(\wb_counter[13] ),
    .A2(_02061_),
    .Z(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07383_ (.A1(net60),
    .A2(_02059_),
    .B(_02065_),
    .ZN(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07384_ (.A1(_02056_),
    .A2(_02067_),
    .B(_02068_),
    .ZN(_00097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07385_ (.A1(_01894_),
    .A2(_02061_),
    .ZN(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07386_ (.A1(_01901_),
    .A2(_02069_),
    .Z(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07387_ (.A1(net61),
    .A2(_02059_),
    .B(_02065_),
    .ZN(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07388_ (.A1(_02056_),
    .A2(_02070_),
    .B(_02071_),
    .ZN(_00098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07389_ (.I(_02012_),
    .Z(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07390_ (.I(_02072_),
    .Z(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07391_ (.A1(\wb_counter[14] ),
    .A2(\wb_counter[15] ),
    .A3(_02069_),
    .ZN(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07392_ (.A1(\wb_counter[14] ),
    .A2(_02069_),
    .ZN(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07393_ (.A1(_01907_),
    .A2(_02075_),
    .ZN(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07394_ (.A1(_02074_),
    .A2(_02076_),
    .ZN(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07395_ (.I(_02026_),
    .Z(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07396_ (.A1(net62),
    .A2(_02078_),
    .B(_02065_),
    .ZN(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07397_ (.A1(_02073_),
    .A2(_02077_),
    .B(_02079_),
    .ZN(_00099_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07398_ (.A1(\wb_counter[16] ),
    .A2(_02074_),
    .Z(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07399_ (.I(_01751_),
    .Z(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07400_ (.I(_02081_),
    .Z(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07401_ (.A1(net63),
    .A2(_02078_),
    .B(_02082_),
    .ZN(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07402_ (.A1(_02073_),
    .A2(_02080_),
    .B(_02083_),
    .ZN(_00100_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07403_ (.I(\wb_counter[16] ),
    .ZN(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07404_ (.A1(_02084_),
    .A2(_02074_),
    .ZN(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07405_ (.A1(\wb_counter[17] ),
    .A2(_02085_),
    .ZN(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07406_ (.A1(net64),
    .A2(_02078_),
    .B(_02082_),
    .ZN(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07407_ (.A1(_02073_),
    .A2(_02086_),
    .B(_02087_),
    .ZN(_00101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07408_ (.A1(\wb_counter[17] ),
    .A2(_02085_),
    .ZN(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07409_ (.A1(\wb_counter[18] ),
    .A2(_02088_),
    .Z(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07410_ (.A1(net351),
    .A2(_02078_),
    .B(_02082_),
    .ZN(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07411_ (.A1(_02073_),
    .A2(_02089_),
    .B(_02090_),
    .ZN(_00102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07412_ (.I(_02072_),
    .Z(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07413_ (.A1(\wb_counter[17] ),
    .A2(\wb_counter[18] ),
    .A3(_02085_),
    .ZN(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07414_ (.A1(\wb_counter[19] ),
    .A2(_02092_),
    .Z(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07415_ (.I(_02022_),
    .Z(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07416_ (.A1(net66),
    .A2(_02094_),
    .B(_02082_),
    .ZN(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07417_ (.A1(_02091_),
    .A2(_02093_),
    .B(_02095_),
    .ZN(_00103_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07418_ (.I(\wb_counter[19] ),
    .ZN(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07419_ (.A1(_02096_),
    .A2(_02092_),
    .ZN(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07420_ (.A1(\wb_counter[20] ),
    .A2(_02097_),
    .ZN(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07421_ (.I(_02081_),
    .Z(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07422_ (.A1(net68),
    .A2(_02094_),
    .B(_02099_),
    .ZN(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07423_ (.A1(_02091_),
    .A2(_02098_),
    .B(_02100_),
    .ZN(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07424_ (.A1(\wb_counter[20] ),
    .A2(_02097_),
    .ZN(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07425_ (.A1(\wb_counter[21] ),
    .A2(_02101_),
    .Z(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07426_ (.A1(net69),
    .A2(_02094_),
    .B(_02099_),
    .ZN(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07427_ (.A1(_02091_),
    .A2(_02102_),
    .B(_02103_),
    .ZN(_00105_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07428_ (.A1(\wb_counter[20] ),
    .A2(\wb_counter[21] ),
    .A3(_02097_),
    .ZN(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07429_ (.A1(\wb_counter[22] ),
    .A2(_02104_),
    .Z(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07430_ (.A1(net70),
    .A2(_02094_),
    .B(_02099_),
    .ZN(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07431_ (.A1(_02091_),
    .A2(_02105_),
    .B(_02106_),
    .ZN(_00106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07432_ (.I(_02072_),
    .Z(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07433_ (.I(\wb_counter[22] ),
    .ZN(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07434_ (.A1(_02108_),
    .A2(_02104_),
    .ZN(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07435_ (.A1(\wb_counter[23] ),
    .A2(_02109_),
    .ZN(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07436_ (.I(_02022_),
    .Z(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07437_ (.A1(net71),
    .A2(_02111_),
    .B(_02099_),
    .ZN(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07438_ (.A1(_02107_),
    .A2(_02110_),
    .B(_02112_),
    .ZN(_00107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07439_ (.A1(\wb_counter[23] ),
    .A2(_02109_),
    .ZN(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07440_ (.A1(\wb_counter[24] ),
    .A2(_02113_),
    .Z(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07441_ (.I(_02081_),
    .Z(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07442_ (.A1(net72),
    .A2(_02111_),
    .B(_02115_),
    .ZN(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07443_ (.A1(_02107_),
    .A2(_02114_),
    .B(_02116_),
    .ZN(_00108_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07444_ (.A1(\wb_counter[23] ),
    .A2(\wb_counter[24] ),
    .A3(_02109_),
    .ZN(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07445_ (.A1(\wb_counter[25] ),
    .A2(_02117_),
    .Z(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07446_ (.A1(net73),
    .A2(_02111_),
    .B(_02115_),
    .ZN(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07447_ (.A1(_02107_),
    .A2(_02118_),
    .B(_02119_),
    .ZN(_00109_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07448_ (.I(\wb_counter[25] ),
    .ZN(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07449_ (.A1(_02120_),
    .A2(_02117_),
    .ZN(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07450_ (.A1(\wb_counter[26] ),
    .A2(_02121_),
    .ZN(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07451_ (.A1(net74),
    .A2(_02111_),
    .B(_02115_),
    .ZN(_02123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07452_ (.A1(_02107_),
    .A2(_02122_),
    .B(_02123_),
    .ZN(_00110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07453_ (.I(_02072_),
    .Z(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07454_ (.A1(\wb_counter[26] ),
    .A2(_02121_),
    .ZN(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07455_ (.A1(\wb_counter[27] ),
    .A2(_02125_),
    .Z(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07456_ (.I(_02022_),
    .Z(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07457_ (.A1(net75),
    .A2(_02127_),
    .B(_02115_),
    .ZN(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07458_ (.A1(_02124_),
    .A2(_02126_),
    .B(_02128_),
    .ZN(_00111_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07459_ (.A1(\wb_counter[26] ),
    .A2(\wb_counter[27] ),
    .A3(_02121_),
    .ZN(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07460_ (.A1(\wb_counter[28] ),
    .A2(_02129_),
    .Z(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07461_ (.I(_02081_),
    .Z(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07462_ (.A1(net76),
    .A2(_02127_),
    .B(_02131_),
    .ZN(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07463_ (.A1(_02124_),
    .A2(_02130_),
    .B(_02132_),
    .ZN(_00112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07464_ (.I(\wb_counter[28] ),
    .ZN(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07465_ (.A1(_02133_),
    .A2(_02129_),
    .ZN(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07466_ (.A1(\wb_counter[29] ),
    .A2(_02134_),
    .ZN(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07467_ (.A1(net77),
    .A2(_02127_),
    .B(_02131_),
    .ZN(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07468_ (.A1(_02124_),
    .A2(_02135_),
    .B(_02136_),
    .ZN(_00113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07469_ (.A1(\wb_counter[29] ),
    .A2(_02134_),
    .ZN(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07470_ (.A1(\wb_counter[30] ),
    .A2(_02137_),
    .Z(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07471_ (.A1(net79),
    .A2(_02127_),
    .B(_02131_),
    .ZN(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07472_ (.A1(_02124_),
    .A2(_02138_),
    .B(_02139_),
    .ZN(_00114_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07473_ (.A1(\wb_counter[29] ),
    .A2(\wb_counter[30] ),
    .A3(_02134_),
    .ZN(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07474_ (.A1(\wb_counter[31] ),
    .A2(_02140_),
    .Z(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07475_ (.A1(net80),
    .A2(_02023_),
    .B(_02131_),
    .ZN(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07476_ (.A1(_02014_),
    .A2(_02141_),
    .B(_02142_),
    .ZN(_00115_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07477_ (.I(_00654_),
    .Z(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07478_ (.A1(_02143_),
    .A2(_00645_),
    .A3(_01243_),
    .ZN(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _07479_ (.A1(_01408_),
    .A2(_01366_),
    .ZN(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07480_ (.A1(_02145_),
    .A2(_01676_),
    .ZN(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07481_ (.A1(_01661_),
    .A2(_02146_),
    .Z(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07482_ (.A1(_01663_),
    .A2(_02147_),
    .ZN(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07483_ (.I(_00957_),
    .Z(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07484_ (.A1(_01228_),
    .A2(_01673_),
    .B(_02145_),
    .ZN(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07485_ (.A1(_02149_),
    .A2(_02150_),
    .ZN(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07486_ (.I(_02143_),
    .Z(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07487_ (.I(_00651_),
    .Z(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07488_ (.A1(_02152_),
    .A2(_02153_),
    .ZN(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07489_ (.A1(_02144_),
    .A2(_02148_),
    .B(_02151_),
    .C(_02154_),
    .ZN(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07490_ (.A1(_01469_),
    .A2(_01408_),
    .ZN(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07491_ (.I(_01508_),
    .Z(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07492_ (.I(_02157_),
    .Z(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07493_ (.A1(_01407_),
    .A2(_01390_),
    .ZN(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07494_ (.I(_02159_),
    .Z(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07495_ (.I(_02160_),
    .Z(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07496_ (.I(_00911_),
    .Z(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07497_ (.A1(_01362_),
    .A2(_02159_),
    .ZN(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07498_ (.A1(_02162_),
    .A2(_02161_),
    .B1(_02163_),
    .B2(_00921_),
    .ZN(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _07499_ (.A1(_02158_),
    .A2(_00906_),
    .A3(_02161_),
    .B(_02164_),
    .ZN(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _07500_ (.A1(_01378_),
    .A2(_01403_),
    .ZN(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07501_ (.A1(_01508_),
    .A2(_02166_),
    .ZN(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07502_ (.I(_02167_),
    .Z(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07503_ (.A1(_00920_),
    .A2(_00979_),
    .Z(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07504_ (.A1(_02157_),
    .A2(_02160_),
    .ZN(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07505_ (.I(_02170_),
    .Z(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07506_ (.A1(_00985_),
    .A2(_02171_),
    .ZN(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _07507_ (.A1(_01633_),
    .A2(_02166_),
    .B1(_02168_),
    .B2(_02169_),
    .C(_02172_),
    .ZN(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07508_ (.A1(_01084_),
    .A2(_01085_),
    .A3(_02168_),
    .ZN(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _07509_ (.A1(_01086_),
    .A2(_02161_),
    .B1(_02171_),
    .B2(_01619_),
    .C(_02174_),
    .ZN(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07510_ (.A1(_01588_),
    .A2(_01047_),
    .B(_01067_),
    .ZN(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07511_ (.A1(_02176_),
    .A2(_02168_),
    .ZN(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _07512_ (.A1(_01588_),
    .A2(_02160_),
    .B1(_02171_),
    .B2(_01074_),
    .C(_02177_),
    .ZN(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07513_ (.A1(_01099_),
    .A2(_02168_),
    .ZN(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _07514_ (.A1(_01601_),
    .A2(_02161_),
    .B1(_02171_),
    .B2(_01098_),
    .C(_02179_),
    .ZN(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _07515_ (.A1(_01047_),
    .A2(_01050_),
    .A3(_02167_),
    .Z(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07516_ (.A1(_01053_),
    .A2(_01054_),
    .ZN(_02182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07517_ (.A1(_01574_),
    .A2(_02160_),
    .B1(_02170_),
    .B2(_02182_),
    .ZN(_02183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07518_ (.A1(_02181_),
    .A2(_02183_),
    .ZN(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07519_ (.I(_00973_),
    .Z(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07520_ (.A1(_02185_),
    .A2(_02166_),
    .Z(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07521_ (.I(_01005_),
    .Z(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07522_ (.A1(_02187_),
    .A2(_02159_),
    .B(_02163_),
    .ZN(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07523_ (.A1(_01024_),
    .A2(_02188_),
    .ZN(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07524_ (.A1(_02184_),
    .A2(_02186_),
    .A3(_02189_),
    .ZN(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07525_ (.A1(_02175_),
    .A2(_02178_),
    .A3(_02180_),
    .A4(_02190_),
    .ZN(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07526_ (.A1(_02165_),
    .A2(_02173_),
    .A3(_02191_),
    .ZN(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07527_ (.A1(_02156_),
    .A2(_02192_),
    .ZN(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07528_ (.A1(\as2650.debug_psl[6] ),
    .A2(_00785_),
    .Z(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07529_ (.A1(\as2650.debug_psl[7] ),
    .A2(_00803_),
    .Z(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07530_ (.A1(_02194_),
    .A2(_02195_),
    .ZN(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07531_ (.A1(_01507_),
    .A2(_02196_),
    .ZN(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07532_ (.A1(_01443_),
    .A2(_02156_),
    .A3(_02197_),
    .ZN(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07533_ (.A1(_01461_),
    .A2(_01379_),
    .ZN(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07534_ (.A1(_01441_),
    .A2(_02199_),
    .ZN(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07535_ (.A1(_00713_),
    .A2(_00717_),
    .ZN(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07536_ (.A1(_02201_),
    .A2(_01506_),
    .ZN(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07537_ (.A1(_01400_),
    .A2(_02200_),
    .A3(_02202_),
    .ZN(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07538_ (.I(_02203_),
    .Z(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07539_ (.I(_02204_),
    .Z(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07540_ (.I(_00687_),
    .Z(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _07541_ (.A1(_02206_),
    .A2(_00722_),
    .A3(_01506_),
    .A4(_01659_),
    .ZN(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07542_ (.A1(_02196_),
    .A2(_02200_),
    .B(_02207_),
    .C(_01179_),
    .ZN(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07543_ (.A1(_02198_),
    .A2(_02205_),
    .A3(_02208_),
    .ZN(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07544_ (.A1(_02193_),
    .A2(_02209_),
    .ZN(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07545_ (.I(_01403_),
    .Z(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07546_ (.I(_01379_),
    .Z(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07547_ (.A1(_02212_),
    .A2(_01365_),
    .ZN(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07548_ (.A1(_02143_),
    .A2(_02153_),
    .B1(_02211_),
    .B2(_02213_),
    .ZN(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07549_ (.I(_02214_),
    .ZN(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07550_ (.A1(_02210_),
    .A2(_02215_),
    .ZN(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07551_ (.A1(_01346_),
    .A2(_01351_),
    .A3(_02216_),
    .ZN(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _07552_ (.A1(_02217_),
    .A2(_02155_),
    .Z(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07553_ (.I(_02218_),
    .ZN(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07554_ (.I(_02219_),
    .Z(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07555_ (.I(_02220_),
    .Z(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07556_ (.I(\as2650.PC[0] ),
    .Z(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07557_ (.I(_00955_),
    .Z(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07558_ (.A1(_02222_),
    .A2(_02223_),
    .Z(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07559_ (.I(\as2650.debug_psl[0] ),
    .Z(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07560_ (.I(_02225_),
    .Z(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07561_ (.I(_02226_),
    .Z(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07562_ (.I(_01505_),
    .Z(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07563_ (.I(_02228_),
    .Z(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07564_ (.I(_01511_),
    .Z(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _07565_ (.A1(_01618_),
    .A2(_02230_),
    .Z(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07566_ (.A1(_01514_),
    .A2(_01344_),
    .A3(_01350_),
    .ZN(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07567_ (.I(_02232_),
    .Z(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07568_ (.I(_02233_),
    .Z(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07569_ (.I(_02234_),
    .Z(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07570_ (.A1(_02229_),
    .A2(_02231_),
    .A3(_02235_),
    .ZN(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07571_ (.I(_02236_),
    .Z(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07572_ (.I(_02237_),
    .Z(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07573_ (.I(_01320_),
    .Z(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07574_ (.I(_02236_),
    .Z(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07575_ (.I(_02240_),
    .Z(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07576_ (.A1(_02239_),
    .A2(_02241_),
    .ZN(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07577_ (.A1(_02227_),
    .A2(_02238_),
    .B(_02242_),
    .C(_02220_),
    .ZN(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07578_ (.A1(_02221_),
    .A2(_02224_),
    .B(_02243_),
    .ZN(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07579_ (.I(_02244_),
    .Z(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _07580_ (.I(\as2650.debug_psu[2] ),
    .ZN(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07581_ (.I(_02246_),
    .Z(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07582_ (.I(_01880_),
    .Z(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07583_ (.A1(_01847_),
    .A2(_01858_),
    .Z(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07584_ (.I(_02249_),
    .Z(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07585_ (.I(_02250_),
    .Z(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07586_ (.I(_02251_),
    .Z(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07587_ (.I(_02252_),
    .Z(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07588_ (.I(_02253_),
    .Z(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07589_ (.I(_02254_),
    .Z(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07590_ (.I(_02230_),
    .Z(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07591_ (.A1(_01618_),
    .A2(_02256_),
    .ZN(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07592_ (.I(_00677_),
    .Z(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07593_ (.A1(_02258_),
    .A2(_01654_),
    .A3(_01429_),
    .ZN(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07594_ (.I(_02259_),
    .Z(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07595_ (.I(_02260_),
    .Z(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07596_ (.A1(_02257_),
    .A2(_02261_),
    .B(_02219_),
    .ZN(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07597_ (.I(_02262_),
    .Z(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07598_ (.I(_02263_),
    .Z(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _07599_ (.A1(_02247_),
    .A2(_02248_),
    .A3(_02255_),
    .A4(_02264_),
    .ZN(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07600_ (.I(_02265_),
    .Z(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07601_ (.I0(_02245_),
    .I1(\as2650.stack[11][0] ),
    .S(_02266_),
    .Z(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07602_ (.I(_02267_),
    .Z(_00117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07603_ (.I(\as2650.debug_psl[1] ),
    .Z(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07604_ (.I(_02268_),
    .Z(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07605_ (.I(_02237_),
    .Z(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07606_ (.I(_02240_),
    .Z(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07607_ (.A1(_01564_),
    .A2(_02271_),
    .ZN(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07608_ (.I(_02220_),
    .Z(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07609_ (.A1(_02269_),
    .A2(_02270_),
    .B(_02272_),
    .C(_02273_),
    .ZN(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07610_ (.I(\as2650.PC[1] ),
    .Z(_02275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07611_ (.I(_02275_),
    .Z(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07612_ (.I(_00659_),
    .Z(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07613_ (.I(_02277_),
    .Z(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07614_ (.I(_02218_),
    .Z(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07615_ (.I(_02277_),
    .Z(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07616_ (.I(_00951_),
    .Z(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07617_ (.A1(_02281_),
    .A2(_02276_),
    .Z(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07618_ (.I(_02282_),
    .Z(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07619_ (.A1(_02280_),
    .A2(_02283_),
    .ZN(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07620_ (.A1(_02276_),
    .A2(_02278_),
    .B(_02279_),
    .C(_02284_),
    .ZN(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07621_ (.A1(_02274_),
    .A2(_02285_),
    .ZN(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07622_ (.I(_02286_),
    .Z(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07623_ (.I0(_02287_),
    .I1(\as2650.stack[11][1] ),
    .S(_02266_),
    .Z(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07624_ (.I(_02288_),
    .Z(_00118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07625_ (.I(\as2650.debug_psl[2] ),
    .Z(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07626_ (.I(_02237_),
    .Z(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07627_ (.I(_01333_),
    .Z(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07628_ (.I(_02240_),
    .Z(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07629_ (.A1(_02291_),
    .A2(_02292_),
    .ZN(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07630_ (.A1(_02289_),
    .A2(_02290_),
    .B(_02293_),
    .C(_02273_),
    .ZN(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07631_ (.I(\as2650.PC[2] ),
    .Z(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07632_ (.I(_02295_),
    .Z(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07633_ (.A1(\as2650.PC[0] ),
    .A2(_02275_),
    .ZN(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07634_ (.A1(_02295_),
    .A2(_02297_),
    .Z(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07635_ (.A1(_02280_),
    .A2(_02298_),
    .ZN(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07636_ (.A1(_02296_),
    .A2(_02278_),
    .B(_02279_),
    .C(_02299_),
    .ZN(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07637_ (.A1(_02294_),
    .A2(_02300_),
    .ZN(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07638_ (.I(_02301_),
    .Z(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07639_ (.I0(_02302_),
    .I1(\as2650.stack[11][2] ),
    .S(_02266_),
    .Z(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07640_ (.I(_02303_),
    .Z(_00119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07641_ (.A1(_01592_),
    .A2(_02292_),
    .ZN(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07642_ (.A1(_01804_),
    .A2(_02290_),
    .B(_02304_),
    .C(_02273_),
    .ZN(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07643_ (.I(\as2650.PC[3] ),
    .Z(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07644_ (.I(_02218_),
    .Z(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07645_ (.I(_02307_),
    .Z(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07646_ (.A1(\as2650.PC[0] ),
    .A2(_02275_),
    .A3(\as2650.PC[2] ),
    .ZN(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07647_ (.A1(_02306_),
    .A2(_02309_),
    .Z(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07648_ (.I(_02310_),
    .Z(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07649_ (.A1(_02280_),
    .A2(_02311_),
    .ZN(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07650_ (.A1(_02306_),
    .A2(_02278_),
    .B(_02308_),
    .C(_02312_),
    .ZN(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07651_ (.A1(_02305_),
    .A2(_02313_),
    .ZN(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07652_ (.I(_02314_),
    .Z(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07653_ (.I0(_02315_),
    .I1(\as2650.stack[11][3] ),
    .S(_02266_),
    .Z(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07654_ (.I(_02316_),
    .Z(_00120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07655_ (.I(_00634_),
    .Z(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07656_ (.A1(_02317_),
    .A2(_02292_),
    .ZN(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07657_ (.I(_02219_),
    .Z(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07658_ (.A1(_01814_),
    .A2(_02290_),
    .B(_02318_),
    .C(_02319_),
    .ZN(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07659_ (.I(\as2650.PC[4] ),
    .Z(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07660_ (.I(_02321_),
    .Z(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07661_ (.A1(_00946_),
    .A2(_02309_),
    .ZN(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _07662_ (.A1(_02321_),
    .A2(_02323_),
    .ZN(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07663_ (.A1(_02280_),
    .A2(_02324_),
    .ZN(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07664_ (.A1(_02322_),
    .A2(_02278_),
    .B(_02308_),
    .C(_02325_),
    .ZN(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07665_ (.A1(_02320_),
    .A2(_02326_),
    .ZN(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07666_ (.I(_02327_),
    .Z(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07667_ (.I(_02265_),
    .Z(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07668_ (.I0(_02328_),
    .I1(\as2650.stack[11][4] ),
    .S(_02329_),
    .Z(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07669_ (.I(_02330_),
    .Z(_00121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07670_ (.I(_01622_),
    .Z(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07671_ (.A1(_02331_),
    .A2(_02292_),
    .ZN(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07672_ (.A1(_01827_),
    .A2(_02290_),
    .B(_02332_),
    .C(_02319_),
    .ZN(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07673_ (.I(\as2650.PC[5] ),
    .Z(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07674_ (.I(_02334_),
    .Z(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07675_ (.I(_02277_),
    .Z(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _07676_ (.A1(\as2650.PC[4] ),
    .A2(_02323_),
    .Z(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07677_ (.A1(_02335_),
    .A2(_02337_),
    .ZN(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07678_ (.A1(_02277_),
    .A2(_02338_),
    .ZN(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07679_ (.A1(_02335_),
    .A2(_02336_),
    .B(_02308_),
    .C(_02339_),
    .ZN(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07680_ (.A1(_02333_),
    .A2(_02340_),
    .ZN(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07681_ (.I(_02341_),
    .Z(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07682_ (.I0(_02342_),
    .I1(\as2650.stack[11][5] ),
    .S(_02329_),
    .Z(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07683_ (.I(_02343_),
    .Z(_00122_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07684_ (.I(_02237_),
    .Z(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07685_ (.I(_00621_),
    .ZN(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07686_ (.I(_02345_),
    .Z(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07687_ (.I(_02240_),
    .Z(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07688_ (.A1(_02346_),
    .A2(_02347_),
    .ZN(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07689_ (.A1(_01460_),
    .A2(_02344_),
    .B(_02348_),
    .C(_02319_),
    .ZN(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07690_ (.I(\as2650.PC[6] ),
    .Z(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07691_ (.I(_02350_),
    .Z(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07692_ (.A1(\as2650.PC[5] ),
    .A2(_02337_),
    .ZN(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07693_ (.A1(_02350_),
    .A2(_02352_),
    .ZN(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07694_ (.I(_02353_),
    .Z(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07695_ (.A1(_02223_),
    .A2(_02354_),
    .Z(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07696_ (.A1(_02351_),
    .A2(_02336_),
    .B(_02308_),
    .C(_02355_),
    .ZN(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07697_ (.A1(_02349_),
    .A2(_02356_),
    .ZN(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07698_ (.I(_02357_),
    .Z(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07699_ (.I0(_02358_),
    .I1(\as2650.stack[11][6] ),
    .S(_02329_),
    .Z(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07700_ (.I(_02359_),
    .Z(_00123_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07701_ (.I(_01644_),
    .Z(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07702_ (.A1(_02360_),
    .A2(_02347_),
    .ZN(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07703_ (.A1(_01468_),
    .A2(_02344_),
    .B(_02361_),
    .C(_02319_),
    .ZN(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07704_ (.I(_00955_),
    .Z(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07705_ (.I(\as2650.PC[7] ),
    .Z(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07706_ (.I(_02364_),
    .ZN(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07707_ (.A1(_02334_),
    .A2(_02350_),
    .A3(_02337_),
    .ZN(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _07708_ (.A1(_02365_),
    .A2(_02366_),
    .Z(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07709_ (.I(_02367_),
    .Z(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07710_ (.I(_00955_),
    .Z(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07711_ (.A1(_02365_),
    .A2(_02369_),
    .ZN(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07712_ (.I(_02307_),
    .Z(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07713_ (.A1(_02363_),
    .A2(_02368_),
    .B(_02370_),
    .C(_02371_),
    .ZN(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07714_ (.A1(_02362_),
    .A2(_02372_),
    .ZN(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07715_ (.I(_02373_),
    .Z(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07716_ (.I0(_02374_),
    .I1(\as2650.stack[11][7] ),
    .S(_02329_),
    .Z(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07717_ (.I(_02375_),
    .Z(_00124_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07718_ (.I(_00607_),
    .ZN(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07719_ (.A1(_02376_),
    .A2(_02347_),
    .ZN(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07720_ (.I(_02219_),
    .Z(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07721_ (.A1(_01848_),
    .A2(_02344_),
    .B(_02377_),
    .C(_02378_),
    .ZN(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07722_ (.I(\as2650.PC[8] ),
    .Z(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07723_ (.A1(_02365_),
    .A2(_02366_),
    .ZN(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07724_ (.A1(_02380_),
    .A2(_02381_),
    .Z(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07725_ (.I(_02382_),
    .Z(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07726_ (.I(_02383_),
    .Z(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07727_ (.I(_02380_),
    .Z(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07728_ (.I(_02385_),
    .ZN(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07729_ (.A1(_02386_),
    .A2(_02369_),
    .ZN(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07730_ (.A1(_02363_),
    .A2(_02384_),
    .B(_02387_),
    .C(_02279_),
    .ZN(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07731_ (.A1(_02379_),
    .A2(_02388_),
    .ZN(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07732_ (.I(_02389_),
    .Z(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07733_ (.I(_02265_),
    .Z(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07734_ (.I0(_02390_),
    .I1(\as2650.stack[11][8] ),
    .S(_02391_),
    .Z(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07735_ (.I(_02392_),
    .Z(_00125_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _07736_ (.I(_00604_),
    .ZN(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07737_ (.A1(_02393_),
    .A2(_02347_),
    .ZN(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07738_ (.A1(_01860_),
    .A2(_02344_),
    .B(_02394_),
    .C(_02378_),
    .ZN(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07739_ (.I(\as2650.PC[9] ),
    .Z(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07740_ (.A1(_02380_),
    .A2(_02381_),
    .ZN(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _07741_ (.A1(\as2650.PC[9] ),
    .A2(_02397_),
    .ZN(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07742_ (.I(_02398_),
    .Z(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07743_ (.A1(_02223_),
    .A2(_02399_),
    .Z(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07744_ (.A1(_02396_),
    .A2(_02336_),
    .B(_02307_),
    .C(_02400_),
    .ZN(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07745_ (.A1(_02395_),
    .A2(_02401_),
    .ZN(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07746_ (.I(_02402_),
    .Z(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07747_ (.I0(_02403_),
    .I1(\as2650.stack[11][9] ),
    .S(_02391_),
    .Z(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07748_ (.I(_02404_),
    .Z(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07749_ (.I(_01867_),
    .Z(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _07750_ (.I(net172),
    .ZN(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07751_ (.A1(_02406_),
    .A2(_02241_),
    .ZN(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07752_ (.A1(_02405_),
    .A2(_02238_),
    .B(_02407_),
    .C(_02378_),
    .ZN(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07753_ (.I(\as2650.PC[10] ),
    .ZN(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07754_ (.I(_02409_),
    .Z(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07755_ (.A1(_02380_),
    .A2(_02396_),
    .A3(_02381_),
    .ZN(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07756_ (.A1(_02410_),
    .A2(_02411_),
    .Z(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07757_ (.I(_02412_),
    .Z(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07758_ (.A1(_02410_),
    .A2(_02369_),
    .ZN(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07759_ (.A1(_02363_),
    .A2(_02413_),
    .B(_02414_),
    .C(_02279_),
    .ZN(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07760_ (.A1(_02408_),
    .A2(_02415_),
    .ZN(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07761_ (.I(_02416_),
    .Z(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07762_ (.I0(_02417_),
    .I1(\as2650.stack[11][10] ),
    .S(_02391_),
    .Z(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07763_ (.I(_02418_),
    .Z(_00127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07764_ (.I(\as2650.PC[11] ),
    .Z(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07765_ (.A1(_02409_),
    .A2(_02411_),
    .ZN(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07766_ (.A1(_02419_),
    .A2(_02420_),
    .Z(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07767_ (.I(_02421_),
    .Z(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07768_ (.I(_02419_),
    .ZN(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07769_ (.A1(_02423_),
    .A2(_02369_),
    .ZN(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07770_ (.A1(_02363_),
    .A2(_02422_),
    .B(_02424_),
    .ZN(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07771_ (.I(_01879_),
    .Z(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07772_ (.I(net173),
    .ZN(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07773_ (.A1(_02427_),
    .A2(_02241_),
    .ZN(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07774_ (.A1(_02426_),
    .A2(_02238_),
    .B(_02428_),
    .C(_02220_),
    .ZN(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07775_ (.A1(_02221_),
    .A2(_02425_),
    .B(_02429_),
    .ZN(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07776_ (.I(_02430_),
    .Z(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07777_ (.I0(_02431_),
    .I1(\as2650.stack[11][11] ),
    .S(_02391_),
    .Z(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07778_ (.I(_02432_),
    .Z(_00128_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07779_ (.I(_00594_),
    .ZN(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07780_ (.I(_02433_),
    .Z(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07781_ (.A1(_02434_),
    .A2(_02241_),
    .ZN(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07782_ (.A1(_01888_),
    .A2(_02238_),
    .B(_02435_),
    .C(_02378_),
    .ZN(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07783_ (.I(\as2650.PC[12] ),
    .Z(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07784_ (.A1(_02419_),
    .A2(_02420_),
    .ZN(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07785_ (.I(_02438_),
    .ZN(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07786_ (.A1(_02437_),
    .A2(_02439_),
    .Z(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07787_ (.I(_02440_),
    .Z(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07788_ (.A1(_02223_),
    .A2(_02441_),
    .Z(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07789_ (.A1(_02437_),
    .A2(_02336_),
    .B(_02307_),
    .C(_02442_),
    .ZN(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07790_ (.A1(_02436_),
    .A2(_02443_),
    .ZN(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07791_ (.I(_02444_),
    .Z(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07792_ (.I(_02265_),
    .Z(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07793_ (.I0(_02445_),
    .I1(\as2650.stack[11][12] ),
    .S(_02446_),
    .Z(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07794_ (.I(_02447_),
    .Z(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07795_ (.I(\as2650.page_reg[0] ),
    .Z(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07796_ (.A1(_02448_),
    .A2(_02371_),
    .ZN(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07797_ (.I(_00591_),
    .ZN(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07798_ (.I(_02450_),
    .Z(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07799_ (.A1(_02451_),
    .A2(_02271_),
    .ZN(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07800_ (.A1(_01897_),
    .A2(_02270_),
    .B(_02452_),
    .C(_02221_),
    .ZN(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07801_ (.A1(_02449_),
    .A2(_02453_),
    .ZN(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07802_ (.I(_02454_),
    .Z(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07803_ (.I0(_02455_),
    .I1(\as2650.stack[11][13] ),
    .S(_02446_),
    .Z(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07804_ (.I(_02456_),
    .Z(_00130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07805_ (.I(\as2650.page_reg[1] ),
    .Z(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07806_ (.A1(_02457_),
    .A2(_02371_),
    .ZN(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07807_ (.I(_00589_),
    .Z(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _07808_ (.I(_02459_),
    .ZN(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07809_ (.A1(_02460_),
    .A2(_02271_),
    .ZN(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07810_ (.A1(net253),
    .A2(_02270_),
    .B(_02461_),
    .C(_02221_),
    .ZN(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07811_ (.A1(_02458_),
    .A2(_02462_),
    .ZN(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07812_ (.I(_02463_),
    .Z(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07813_ (.I0(_02464_),
    .I1(\as2650.stack[11][14] ),
    .S(_02446_),
    .Z(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07814_ (.I(_02465_),
    .Z(_00131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07815_ (.I(\as2650.page_reg[2] ),
    .Z(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07816_ (.A1(_02466_),
    .A2(_02371_),
    .ZN(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07817_ (.I(_00585_),
    .ZN(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07818_ (.I(_02468_),
    .Z(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07819_ (.A1(_02469_),
    .A2(_02271_),
    .ZN(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07820_ (.A1(_01910_),
    .A2(_02270_),
    .B(_02470_),
    .C(_02273_),
    .ZN(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07821_ (.A1(_02467_),
    .A2(_02471_),
    .ZN(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07822_ (.I(_02472_),
    .Z(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07823_ (.I0(_02473_),
    .I1(\as2650.stack[11][15] ),
    .S(_02446_),
    .Z(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07824_ (.I(_02474_),
    .Z(_00132_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07825_ (.I(_01858_),
    .ZN(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07826_ (.A1(_01847_),
    .A2(_02475_),
    .ZN(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07827_ (.I(_02476_),
    .Z(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07828_ (.I(_02477_),
    .Z(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07829_ (.I(_02478_),
    .Z(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07830_ (.I(_02479_),
    .Z(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07831_ (.I(_02480_),
    .Z(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07832_ (.I(_02481_),
    .Z(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07833_ (.I(_02231_),
    .Z(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07834_ (.I(_02234_),
    .Z(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07835_ (.A1(_02483_),
    .A2(_02484_),
    .B(_02218_),
    .ZN(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07836_ (.A1(_01868_),
    .A2(_01880_),
    .A3(_02485_),
    .ZN(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _07837_ (.A1(_02482_),
    .A2(_02486_),
    .ZN(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07838_ (.I(_02487_),
    .Z(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07839_ (.I0(_02245_),
    .I1(\as2650.stack[2][0] ),
    .S(_02488_),
    .Z(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07840_ (.I(_02489_),
    .Z(_00133_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07841_ (.I0(_02287_),
    .I1(\as2650.stack[2][1] ),
    .S(_02488_),
    .Z(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07842_ (.I(_02490_),
    .Z(_00134_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07843_ (.I0(_02302_),
    .I1(\as2650.stack[2][2] ),
    .S(_02488_),
    .Z(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07844_ (.I(_02491_),
    .Z(_00135_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07845_ (.I0(_02315_),
    .I1(\as2650.stack[2][3] ),
    .S(_02488_),
    .Z(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07846_ (.I(_02492_),
    .Z(_00136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07847_ (.I(_02487_),
    .Z(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07848_ (.I0(_02328_),
    .I1(\as2650.stack[2][4] ),
    .S(_02493_),
    .Z(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07849_ (.I(_02494_),
    .Z(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07850_ (.I0(_02342_),
    .I1(\as2650.stack[2][5] ),
    .S(_02493_),
    .Z(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07851_ (.I(_02495_),
    .Z(_00138_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07852_ (.I0(_02358_),
    .I1(\as2650.stack[2][6] ),
    .S(_02493_),
    .Z(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07853_ (.I(_02496_),
    .Z(_00139_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07854_ (.I0(_02374_),
    .I1(\as2650.stack[2][7] ),
    .S(_02493_),
    .Z(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07855_ (.I(_02497_),
    .Z(_00140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07856_ (.I(_02487_),
    .Z(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07857_ (.I0(_02390_),
    .I1(\as2650.stack[2][8] ),
    .S(_02498_),
    .Z(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07858_ (.I(_02499_),
    .Z(_00141_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07859_ (.I0(_02403_),
    .I1(\as2650.stack[2][9] ),
    .S(_02498_),
    .Z(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07860_ (.I(_02500_),
    .Z(_00142_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07861_ (.I0(_02417_),
    .I1(\as2650.stack[2][10] ),
    .S(_02498_),
    .Z(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07862_ (.I(_02501_),
    .Z(_00143_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07863_ (.I0(_02431_),
    .I1(\as2650.stack[2][11] ),
    .S(_02498_),
    .Z(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07864_ (.I(_02502_),
    .Z(_00144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07865_ (.I(_02487_),
    .Z(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07866_ (.I0(_02445_),
    .I1(\as2650.stack[2][12] ),
    .S(_02503_),
    .Z(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07867_ (.I(_02504_),
    .Z(_00145_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07868_ (.I0(_02455_),
    .I1(\as2650.stack[2][13] ),
    .S(_02503_),
    .Z(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07869_ (.I(_02505_),
    .Z(_00146_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07870_ (.I0(_02464_),
    .I1(\as2650.stack[2][14] ),
    .S(_02503_),
    .Z(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07871_ (.I(_02506_),
    .Z(_00147_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07872_ (.I0(_02473_),
    .I1(\as2650.stack[2][15] ),
    .S(_02503_),
    .Z(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07873_ (.I(_02507_),
    .Z(_00148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _07874_ (.A1(_02255_),
    .A2(_02486_),
    .ZN(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07875_ (.I(_02508_),
    .Z(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07876_ (.I0(_02245_),
    .I1(\as2650.stack[3][0] ),
    .S(_02509_),
    .Z(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07877_ (.I(_02510_),
    .Z(_00149_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07878_ (.I0(_02287_),
    .I1(\as2650.stack[3][1] ),
    .S(_02509_),
    .Z(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07879_ (.I(_02511_),
    .Z(_00150_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07880_ (.I0(_02302_),
    .I1(\as2650.stack[3][2] ),
    .S(_02509_),
    .Z(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07881_ (.I(_02512_),
    .Z(_00151_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07882_ (.I0(_02315_),
    .I1(\as2650.stack[3][3] ),
    .S(_02509_),
    .Z(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07883_ (.I(_02513_),
    .Z(_00152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07884_ (.I(_02508_),
    .Z(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07885_ (.I0(_02328_),
    .I1(\as2650.stack[3][4] ),
    .S(_02514_),
    .Z(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07886_ (.I(_02515_),
    .Z(_00153_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07887_ (.I0(_02342_),
    .I1(\as2650.stack[3][5] ),
    .S(_02514_),
    .Z(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07888_ (.I(_02516_),
    .Z(_00154_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07889_ (.I0(_02358_),
    .I1(\as2650.stack[3][6] ),
    .S(_02514_),
    .Z(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07890_ (.I(_02517_),
    .Z(_00155_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07891_ (.I0(_02374_),
    .I1(\as2650.stack[3][7] ),
    .S(_02514_),
    .Z(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07892_ (.I(_02518_),
    .Z(_00156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07893_ (.I(_02508_),
    .Z(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07894_ (.I0(_02390_),
    .I1(\as2650.stack[3][8] ),
    .S(_02519_),
    .Z(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07895_ (.I(_02520_),
    .Z(_00157_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07896_ (.I0(_02403_),
    .I1(\as2650.stack[3][9] ),
    .S(_02519_),
    .Z(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07897_ (.I(_02521_),
    .Z(_00158_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07898_ (.I0(_02417_),
    .I1(\as2650.stack[3][10] ),
    .S(_02519_),
    .Z(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07899_ (.I(_02522_),
    .Z(_00159_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07900_ (.I0(_02431_),
    .I1(\as2650.stack[3][11] ),
    .S(_02519_),
    .Z(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07901_ (.I(_02523_),
    .Z(_00160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07902_ (.I(_02508_),
    .Z(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07903_ (.I0(_02445_),
    .I1(\as2650.stack[3][12] ),
    .S(_02524_),
    .Z(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07904_ (.I(_02525_),
    .Z(_00161_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07905_ (.I0(_02455_),
    .I1(\as2650.stack[3][13] ),
    .S(_02524_),
    .Z(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07906_ (.I(_02526_),
    .Z(_00162_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07907_ (.I0(_02464_),
    .I1(\as2650.stack[3][14] ),
    .S(_02524_),
    .Z(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07908_ (.I(_02527_),
    .Z(_00163_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07909_ (.I0(_02473_),
    .I1(\as2650.stack[3][15] ),
    .S(_02524_),
    .Z(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07910_ (.I(_02528_),
    .Z(_00164_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07911_ (.I(\as2650.debug_psu[3] ),
    .ZN(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07912_ (.I(_02529_),
    .Z(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07913_ (.I(_02530_),
    .Z(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _07914_ (.A1(\as2650.debug_psu[0] ),
    .A2(\as2650.debug_psu[1] ),
    .Z(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _07915_ (.A1(\as2650.debug_psu[2] ),
    .A2(_02532_),
    .ZN(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07916_ (.A1(_02531_),
    .A2(_02264_),
    .A3(_02533_),
    .ZN(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07917_ (.I(_02534_),
    .Z(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07918_ (.I0(_02245_),
    .I1(\as2650.stack[0][0] ),
    .S(_02535_),
    .Z(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07919_ (.I(_02536_),
    .Z(_00165_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07920_ (.I0(_02287_),
    .I1(\as2650.stack[0][1] ),
    .S(_02535_),
    .Z(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07921_ (.I(_02537_),
    .Z(_00166_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07922_ (.I0(_02302_),
    .I1(\as2650.stack[0][2] ),
    .S(_02535_),
    .Z(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07923_ (.I(_02538_),
    .Z(_00167_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07924_ (.I0(_02315_),
    .I1(\as2650.stack[0][3] ),
    .S(_02535_),
    .Z(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07925_ (.I(_02539_),
    .Z(_00168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07926_ (.I(_02534_),
    .Z(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07927_ (.I0(_02328_),
    .I1(\as2650.stack[0][4] ),
    .S(_02540_),
    .Z(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07928_ (.I(_02541_),
    .Z(_00169_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07929_ (.I0(_02342_),
    .I1(\as2650.stack[0][5] ),
    .S(_02540_),
    .Z(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07930_ (.I(_02542_),
    .Z(_00170_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07931_ (.I0(_02358_),
    .I1(\as2650.stack[0][6] ),
    .S(_02540_),
    .Z(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07932_ (.I(_02543_),
    .Z(_00171_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07933_ (.I0(_02374_),
    .I1(\as2650.stack[0][7] ),
    .S(_02540_),
    .Z(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07934_ (.I(_02544_),
    .Z(_00172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07935_ (.I(_02534_),
    .Z(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07936_ (.I0(_02390_),
    .I1(\as2650.stack[0][8] ),
    .S(_02545_),
    .Z(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07937_ (.I(_02546_),
    .Z(_00173_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07938_ (.I0(_02403_),
    .I1(\as2650.stack[0][9] ),
    .S(_02545_),
    .Z(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07939_ (.I(_02547_),
    .Z(_00174_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07940_ (.I0(_02417_),
    .I1(\as2650.stack[0][10] ),
    .S(_02545_),
    .Z(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07941_ (.I(_02548_),
    .Z(_00175_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07942_ (.I0(_02431_),
    .I1(\as2650.stack[0][11] ),
    .S(_02545_),
    .Z(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07943_ (.I(_02549_),
    .Z(_00176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07944_ (.I(_02534_),
    .Z(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07945_ (.I0(_02445_),
    .I1(\as2650.stack[0][12] ),
    .S(_02550_),
    .Z(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07946_ (.I(_02551_),
    .Z(_00177_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07947_ (.I0(_02455_),
    .I1(\as2650.stack[0][13] ),
    .S(_02550_),
    .Z(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07948_ (.I(_02552_),
    .Z(_00178_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07949_ (.I0(_02464_),
    .I1(\as2650.stack[0][14] ),
    .S(_02550_),
    .Z(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07950_ (.I(_02553_),
    .Z(_00179_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07951_ (.I0(_02473_),
    .I1(\as2650.stack[0][15] ),
    .S(_02550_),
    .Z(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07952_ (.I(_02554_),
    .Z(_00180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07953_ (.I(_02244_),
    .Z(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07954_ (.I(_02262_),
    .Z(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__and4_4 _07955_ (.A1(_02405_),
    .A2(_02426_),
    .A3(_02556_),
    .A4(_02482_),
    .Z(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07956_ (.I(_02557_),
    .Z(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07957_ (.I0(\as2650.stack[14][0] ),
    .I1(_02555_),
    .S(_02558_),
    .Z(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07958_ (.I(_02559_),
    .Z(_00181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07959_ (.I(_02286_),
    .Z(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07960_ (.I0(\as2650.stack[14][1] ),
    .I1(_02560_),
    .S(_02558_),
    .Z(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07961_ (.I(_02561_),
    .Z(_00182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07962_ (.I(_02301_),
    .Z(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07963_ (.I0(\as2650.stack[14][2] ),
    .I1(_02562_),
    .S(_02558_),
    .Z(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07964_ (.I(_02563_),
    .Z(_00183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07965_ (.I(_02314_),
    .Z(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07966_ (.I0(\as2650.stack[14][3] ),
    .I1(_02564_),
    .S(_02558_),
    .Z(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07967_ (.I(_02565_),
    .Z(_00184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07968_ (.I(_02327_),
    .Z(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07969_ (.I(_02557_),
    .Z(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07970_ (.I0(\as2650.stack[14][4] ),
    .I1(_02566_),
    .S(_02567_),
    .Z(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07971_ (.I(_02568_),
    .Z(_00185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07972_ (.I(_02341_),
    .Z(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07973_ (.I0(\as2650.stack[14][5] ),
    .I1(_02569_),
    .S(_02567_),
    .Z(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07974_ (.I(_02570_),
    .Z(_00186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07975_ (.I(_02357_),
    .Z(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07976_ (.I0(\as2650.stack[14][6] ),
    .I1(_02571_),
    .S(_02567_),
    .Z(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07977_ (.I(_02572_),
    .Z(_00187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07978_ (.I(_02373_),
    .Z(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07979_ (.I0(\as2650.stack[14][7] ),
    .I1(_02573_),
    .S(_02567_),
    .Z(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07980_ (.I(_02574_),
    .Z(_00188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07981_ (.I(_02389_),
    .Z(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07982_ (.I(_02557_),
    .Z(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07983_ (.I0(\as2650.stack[14][8] ),
    .I1(_02575_),
    .S(_02576_),
    .Z(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07984_ (.I(_02577_),
    .Z(_00189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07985_ (.I(_02402_),
    .Z(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07986_ (.I0(\as2650.stack[14][9] ),
    .I1(_02578_),
    .S(_02576_),
    .Z(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07987_ (.I(_02579_),
    .Z(_00190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07988_ (.I(_02416_),
    .Z(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07989_ (.I0(\as2650.stack[14][10] ),
    .I1(_02580_),
    .S(_02576_),
    .Z(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07990_ (.I(_02581_),
    .Z(_00191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07991_ (.I(_02430_),
    .Z(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07992_ (.I0(\as2650.stack[14][11] ),
    .I1(_02582_),
    .S(_02576_),
    .Z(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07993_ (.I(_02583_),
    .Z(_00192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07994_ (.I(_02444_),
    .Z(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07995_ (.I(_02557_),
    .Z(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07996_ (.I0(\as2650.stack[14][12] ),
    .I1(_02584_),
    .S(_02585_),
    .Z(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07997_ (.I(_02586_),
    .Z(_00193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07998_ (.I(_02454_),
    .Z(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07999_ (.I0(\as2650.stack[14][13] ),
    .I1(_02587_),
    .S(_02585_),
    .Z(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08000_ (.I(_02588_),
    .Z(_00194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08001_ (.I(_02463_),
    .Z(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08002_ (.I0(\as2650.stack[14][14] ),
    .I1(_02589_),
    .S(_02585_),
    .Z(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08003_ (.I(_02590_),
    .Z(_00195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08004_ (.I(_02472_),
    .Z(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08005_ (.I0(\as2650.stack[14][15] ),
    .I1(_02591_),
    .S(_02585_),
    .Z(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08006_ (.I(_02592_),
    .Z(_00196_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08007_ (.A1(\as2650.debug_psu[0] ),
    .A2(_02475_),
    .Z(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08008_ (.I(_02593_),
    .Z(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08009_ (.I(_02594_),
    .Z(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08010_ (.I(_02595_),
    .Z(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08011_ (.I(_02596_),
    .Z(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08012_ (.I(_02597_),
    .Z(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08013_ (.I(_02598_),
    .Z(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__and4_4 _08014_ (.A1(_02405_),
    .A2(_02426_),
    .A3(_02263_),
    .A4(_02599_),
    .Z(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08015_ (.I(_02600_),
    .Z(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08016_ (.I0(\as2650.stack[13][0] ),
    .I1(_02555_),
    .S(_02601_),
    .Z(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08017_ (.I(_02602_),
    .Z(_00197_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08018_ (.I0(\as2650.stack[13][1] ),
    .I1(_02560_),
    .S(_02601_),
    .Z(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08019_ (.I(_02603_),
    .Z(_00198_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08020_ (.I0(\as2650.stack[13][2] ),
    .I1(_02562_),
    .S(_02601_),
    .Z(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08021_ (.I(_02604_),
    .Z(_00199_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08022_ (.I0(\as2650.stack[13][3] ),
    .I1(_02564_),
    .S(_02601_),
    .Z(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08023_ (.I(_02605_),
    .Z(_00200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08024_ (.I(_02600_),
    .Z(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08025_ (.I0(\as2650.stack[13][4] ),
    .I1(_02566_),
    .S(_02606_),
    .Z(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08026_ (.I(_02607_),
    .Z(_00201_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08027_ (.I0(\as2650.stack[13][5] ),
    .I1(_02569_),
    .S(_02606_),
    .Z(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08028_ (.I(_02608_),
    .Z(_00202_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08029_ (.I0(\as2650.stack[13][6] ),
    .I1(_02571_),
    .S(_02606_),
    .Z(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08030_ (.I(_02609_),
    .Z(_00203_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08031_ (.I0(\as2650.stack[13][7] ),
    .I1(_02573_),
    .S(_02606_),
    .Z(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08032_ (.I(_02610_),
    .Z(_00204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08033_ (.I(_02600_),
    .Z(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08034_ (.I0(\as2650.stack[13][8] ),
    .I1(_02575_),
    .S(_02611_),
    .Z(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08035_ (.I(_02612_),
    .Z(_00205_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08036_ (.I0(\as2650.stack[13][9] ),
    .I1(_02578_),
    .S(_02611_),
    .Z(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08037_ (.I(_02613_),
    .Z(_00206_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08038_ (.I0(\as2650.stack[13][10] ),
    .I1(_02580_),
    .S(_02611_),
    .Z(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08039_ (.I(_02614_),
    .Z(_00207_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08040_ (.I0(\as2650.stack[13][11] ),
    .I1(_02582_),
    .S(_02611_),
    .Z(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08041_ (.I(_02615_),
    .Z(_00208_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08042_ (.I(_02600_),
    .Z(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08043_ (.I0(\as2650.stack[13][12] ),
    .I1(_02584_),
    .S(_02616_),
    .Z(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08044_ (.I(_02617_),
    .Z(_00209_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08045_ (.I0(\as2650.stack[13][13] ),
    .I1(_02587_),
    .S(_02616_),
    .Z(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08046_ (.I(_02618_),
    .Z(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08047_ (.I0(\as2650.stack[13][14] ),
    .I1(_02589_),
    .S(_02616_),
    .Z(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08048_ (.I(_02619_),
    .Z(_00211_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08049_ (.I0(\as2650.stack[13][15] ),
    .I1(_02591_),
    .S(_02616_),
    .Z(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08050_ (.I(_02620_),
    .Z(_00212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08051_ (.I(_02244_),
    .Z(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _08052_ (.A1(_02246_),
    .A2(_02530_),
    .A3(_02485_),
    .A4(_02532_),
    .ZN(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08053_ (.I(net248),
    .Z(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08054_ (.I0(\as2650.stack[12][0] ),
    .I1(_02621_),
    .S(_02623_),
    .Z(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08055_ (.I(_02624_),
    .Z(_00213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08056_ (.I(_02286_),
    .Z(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08057_ (.I0(\as2650.stack[12][1] ),
    .I1(_02625_),
    .S(_02623_),
    .Z(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08058_ (.I(_02626_),
    .Z(_00214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08059_ (.I(_02301_),
    .Z(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08060_ (.I0(\as2650.stack[12][2] ),
    .I1(_02627_),
    .S(_02623_),
    .Z(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08061_ (.I(_02628_),
    .Z(_00215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08062_ (.I(_02314_),
    .Z(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08063_ (.I0(\as2650.stack[12][3] ),
    .I1(_02629_),
    .S(_02623_),
    .Z(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08064_ (.I(_02630_),
    .Z(_00216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08065_ (.I(_02327_),
    .Z(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08066_ (.I(net248),
    .Z(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08067_ (.I0(\as2650.stack[12][4] ),
    .I1(_02631_),
    .S(_02632_),
    .Z(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08068_ (.I(_02633_),
    .Z(_00217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08069_ (.I(_02341_),
    .Z(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08070_ (.I0(\as2650.stack[12][5] ),
    .I1(_02634_),
    .S(_02632_),
    .Z(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08071_ (.I(_02635_),
    .Z(_00218_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08072_ (.I(_02357_),
    .Z(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08073_ (.I0(\as2650.stack[12][6] ),
    .I1(_02636_),
    .S(_02632_),
    .Z(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08074_ (.I(_02637_),
    .Z(_00219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08075_ (.I(_02373_),
    .Z(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08076_ (.I0(\as2650.stack[12][7] ),
    .I1(_02638_),
    .S(_02632_),
    .Z(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08077_ (.I(_02639_),
    .Z(_00220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08078_ (.I(_02389_),
    .Z(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08079_ (.I(net248),
    .Z(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08080_ (.I0(\as2650.stack[12][8] ),
    .I1(_02640_),
    .S(_02641_),
    .Z(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08081_ (.I(_02642_),
    .Z(_00221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08082_ (.I(_02402_),
    .Z(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08083_ (.I0(\as2650.stack[12][9] ),
    .I1(_02643_),
    .S(_02641_),
    .Z(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08084_ (.I(_02644_),
    .Z(_00222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08085_ (.I(_02416_),
    .Z(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08086_ (.I0(\as2650.stack[12][10] ),
    .I1(_02645_),
    .S(_02641_),
    .Z(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08087_ (.I(_02646_),
    .Z(_00223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08088_ (.I(_02430_),
    .Z(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08089_ (.I0(\as2650.stack[12][11] ),
    .I1(_02647_),
    .S(_02641_),
    .Z(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08090_ (.I(_02648_),
    .Z(_00224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08091_ (.I(_02444_),
    .Z(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08092_ (.I(net248),
    .Z(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08093_ (.I0(\as2650.stack[12][12] ),
    .I1(_02649_),
    .S(_02650_),
    .Z(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08094_ (.I(_02651_),
    .Z(_00225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08095_ (.I(_02454_),
    .Z(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08096_ (.I0(\as2650.stack[12][13] ),
    .I1(_02652_),
    .S(_02650_),
    .Z(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08097_ (.I(_02653_),
    .Z(_00226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08098_ (.I(_02463_),
    .Z(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08099_ (.I0(\as2650.stack[12][14] ),
    .I1(_02654_),
    .S(_02650_),
    .Z(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08100_ (.I(_02655_),
    .Z(_00227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08101_ (.I(_02472_),
    .Z(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08102_ (.I0(\as2650.stack[12][15] ),
    .I1(_02656_),
    .S(_02650_),
    .Z(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08103_ (.I(_02657_),
    .Z(_00228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08104_ (.I(_02244_),
    .Z(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08105_ (.A1(_01881_),
    .A2(_02264_),
    .A3(_02533_),
    .ZN(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08106_ (.I(_02659_),
    .Z(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08107_ (.I0(_02658_),
    .I1(\as2650.stack[8][0] ),
    .S(_02660_),
    .Z(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08108_ (.I(_02661_),
    .Z(_00229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08109_ (.I(_02286_),
    .Z(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08110_ (.I0(_02662_),
    .I1(\as2650.stack[8][1] ),
    .S(_02660_),
    .Z(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08111_ (.I(_02663_),
    .Z(_00230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08112_ (.I(_02301_),
    .Z(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08113_ (.I0(_02664_),
    .I1(\as2650.stack[8][2] ),
    .S(_02660_),
    .Z(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08114_ (.I(_02665_),
    .Z(_00231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08115_ (.I(_02314_),
    .Z(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08116_ (.I0(_02666_),
    .I1(\as2650.stack[8][3] ),
    .S(_02660_),
    .Z(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08117_ (.I(_02667_),
    .Z(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08118_ (.I(_02327_),
    .Z(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08119_ (.I(_02659_),
    .Z(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08120_ (.I0(_02668_),
    .I1(\as2650.stack[8][4] ),
    .S(_02669_),
    .Z(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08121_ (.I(_02670_),
    .Z(_00233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08122_ (.I(_02341_),
    .Z(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08123_ (.I0(_02671_),
    .I1(\as2650.stack[8][5] ),
    .S(_02669_),
    .Z(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08124_ (.I(_02672_),
    .Z(_00234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08125_ (.I(_02357_),
    .Z(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08126_ (.I0(_02673_),
    .I1(\as2650.stack[8][6] ),
    .S(_02669_),
    .Z(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08127_ (.I(_02674_),
    .Z(_00235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08128_ (.I(_02373_),
    .Z(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08129_ (.I0(_02675_),
    .I1(\as2650.stack[8][7] ),
    .S(_02669_),
    .Z(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08130_ (.I(_02676_),
    .Z(_00236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08131_ (.I(_02389_),
    .Z(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08132_ (.I(_02659_),
    .Z(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08133_ (.I0(_02677_),
    .I1(\as2650.stack[8][8] ),
    .S(_02678_),
    .Z(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08134_ (.I(_02679_),
    .Z(_00237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08135_ (.I(_02402_),
    .Z(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08136_ (.I0(_02680_),
    .I1(\as2650.stack[8][9] ),
    .S(_02678_),
    .Z(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08137_ (.I(_02681_),
    .Z(_00238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08138_ (.I(_02416_),
    .Z(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08139_ (.I0(_02682_),
    .I1(\as2650.stack[8][10] ),
    .S(_02678_),
    .Z(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08140_ (.I(_02683_),
    .Z(_00239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08141_ (.I(_02430_),
    .Z(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08142_ (.I0(_02684_),
    .I1(\as2650.stack[8][11] ),
    .S(_02678_),
    .Z(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08143_ (.I(_02685_),
    .Z(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08144_ (.I(_02444_),
    .Z(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08145_ (.I(_02659_),
    .Z(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08146_ (.I0(_02686_),
    .I1(\as2650.stack[8][12] ),
    .S(_02687_),
    .Z(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08147_ (.I(_02688_),
    .Z(_00241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08148_ (.I(_02454_),
    .Z(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08149_ (.I0(_02689_),
    .I1(\as2650.stack[8][13] ),
    .S(_02687_),
    .Z(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08150_ (.I(_02690_),
    .Z(_00242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08151_ (.I(_02463_),
    .Z(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08152_ (.I0(_02691_),
    .I1(\as2650.stack[8][14] ),
    .S(_02687_),
    .Z(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08153_ (.I(_02692_),
    .Z(_00243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08154_ (.I(_02472_),
    .Z(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08155_ (.I0(_02693_),
    .I1(\as2650.stack[8][15] ),
    .S(_02687_),
    .Z(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08156_ (.I(_02694_),
    .Z(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08157_ (.A1(_01869_),
    .A2(_02531_),
    .A3(_02255_),
    .A4(_02264_),
    .ZN(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08158_ (.I(_02695_),
    .Z(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08159_ (.I0(_02658_),
    .I1(\as2650.stack[7][0] ),
    .S(_02696_),
    .Z(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08160_ (.I(_02697_),
    .Z(_00245_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08161_ (.I0(_02662_),
    .I1(\as2650.stack[7][1] ),
    .S(_02696_),
    .Z(_02698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08162_ (.I(_02698_),
    .Z(_00246_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08163_ (.I0(_02664_),
    .I1(\as2650.stack[7][2] ),
    .S(_02696_),
    .Z(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08164_ (.I(_02699_),
    .Z(_00247_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08165_ (.I0(_02666_),
    .I1(\as2650.stack[7][3] ),
    .S(_02696_),
    .Z(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08166_ (.I(_02700_),
    .Z(_00248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08167_ (.I(_02695_),
    .Z(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08168_ (.I0(_02668_),
    .I1(\as2650.stack[7][4] ),
    .S(_02701_),
    .Z(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08169_ (.I(_02702_),
    .Z(_00249_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08170_ (.I0(_02671_),
    .I1(\as2650.stack[7][5] ),
    .S(_02701_),
    .Z(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08171_ (.I(_02703_),
    .Z(_00250_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08172_ (.I0(_02673_),
    .I1(\as2650.stack[7][6] ),
    .S(_02701_),
    .Z(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08173_ (.I(_02704_),
    .Z(_00251_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08174_ (.I0(_02675_),
    .I1(\as2650.stack[7][7] ),
    .S(_02701_),
    .Z(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08175_ (.I(_02705_),
    .Z(_00252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08176_ (.I(_02695_),
    .Z(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08177_ (.I0(_02677_),
    .I1(\as2650.stack[7][8] ),
    .S(_02706_),
    .Z(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08178_ (.I(_02707_),
    .Z(_00253_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08179_ (.I0(_02680_),
    .I1(\as2650.stack[7][9] ),
    .S(_02706_),
    .Z(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08180_ (.I(_02708_),
    .Z(_00254_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08181_ (.I0(_02682_),
    .I1(\as2650.stack[7][10] ),
    .S(_02706_),
    .Z(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08182_ (.I(_02709_),
    .Z(_00255_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08183_ (.I0(_02684_),
    .I1(\as2650.stack[7][11] ),
    .S(_02706_),
    .Z(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08184_ (.I(_02710_),
    .Z(_00256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08185_ (.I(_02695_),
    .Z(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08186_ (.I0(_02686_),
    .I1(\as2650.stack[7][12] ),
    .S(_02711_),
    .Z(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08187_ (.I(_02712_),
    .Z(_00257_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08188_ (.I0(_02689_),
    .I1(\as2650.stack[7][13] ),
    .S(_02711_),
    .Z(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08189_ (.I(_02713_),
    .Z(_00258_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08190_ (.I0(_02691_),
    .I1(\as2650.stack[7][14] ),
    .S(_02711_),
    .Z(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08191_ (.I(_02714_),
    .Z(_00259_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08192_ (.I0(_02693_),
    .I1(\as2650.stack[7][15] ),
    .S(_02711_),
    .Z(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08193_ (.I(_02715_),
    .Z(_00260_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _08194_ (.A1(_01868_),
    .A2(_02531_),
    .A3(_02263_),
    .A4(_02482_),
    .Z(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08195_ (.I(_02716_),
    .Z(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08196_ (.I0(\as2650.stack[6][0] ),
    .I1(_02621_),
    .S(_02717_),
    .Z(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08197_ (.I(_02718_),
    .Z(_00261_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08198_ (.I0(\as2650.stack[6][1] ),
    .I1(_02625_),
    .S(_02717_),
    .Z(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08199_ (.I(_02719_),
    .Z(_00262_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08200_ (.I0(\as2650.stack[6][2] ),
    .I1(_02627_),
    .S(_02717_),
    .Z(_02720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08201_ (.I(_02720_),
    .Z(_00263_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08202_ (.I0(\as2650.stack[6][3] ),
    .I1(_02629_),
    .S(_02717_),
    .Z(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08203_ (.I(_02721_),
    .Z(_00264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08204_ (.I(_02716_),
    .Z(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08205_ (.I0(\as2650.stack[6][4] ),
    .I1(_02631_),
    .S(_02722_),
    .Z(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08206_ (.I(_02723_),
    .Z(_00265_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08207_ (.I0(\as2650.stack[6][5] ),
    .I1(_02634_),
    .S(_02722_),
    .Z(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08208_ (.I(_02724_),
    .Z(_00266_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08209_ (.I0(\as2650.stack[6][6] ),
    .I1(_02636_),
    .S(_02722_),
    .Z(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08210_ (.I(_02725_),
    .Z(_00267_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08211_ (.I0(\as2650.stack[6][7] ),
    .I1(_02638_),
    .S(_02722_),
    .Z(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08212_ (.I(_02726_),
    .Z(_00268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08213_ (.I(_02716_),
    .Z(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08214_ (.I0(\as2650.stack[6][8] ),
    .I1(_02640_),
    .S(_02727_),
    .Z(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08215_ (.I(_02728_),
    .Z(_00269_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08216_ (.I0(\as2650.stack[6][9] ),
    .I1(_02643_),
    .S(_02727_),
    .Z(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08217_ (.I(_02729_),
    .Z(_00270_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08218_ (.I0(\as2650.stack[6][10] ),
    .I1(_02645_),
    .S(_02727_),
    .Z(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08219_ (.I(_02730_),
    .Z(_00271_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08220_ (.I0(\as2650.stack[6][11] ),
    .I1(_02647_),
    .S(_02727_),
    .Z(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08221_ (.I(_02731_),
    .Z(_00272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08222_ (.I(_02716_),
    .Z(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08223_ (.I0(\as2650.stack[6][12] ),
    .I1(_02649_),
    .S(_02732_),
    .Z(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08224_ (.I(_02733_),
    .Z(_00273_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08225_ (.I0(\as2650.stack[6][13] ),
    .I1(_02652_),
    .S(_02732_),
    .Z(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08226_ (.I(_02734_),
    .Z(_00274_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08227_ (.I0(\as2650.stack[6][14] ),
    .I1(_02654_),
    .S(_02732_),
    .Z(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08228_ (.I(_02735_),
    .Z(_00275_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08229_ (.I0(\as2650.stack[6][15] ),
    .I1(_02656_),
    .S(_02732_),
    .Z(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08230_ (.I(_02736_),
    .Z(_00276_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _08231_ (.A1(_01868_),
    .A2(_02530_),
    .A3(_02263_),
    .A4(_02599_),
    .Z(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08232_ (.I(_02737_),
    .Z(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08233_ (.I0(\as2650.stack[5][0] ),
    .I1(_02621_),
    .S(_02738_),
    .Z(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08234_ (.I(_02739_),
    .Z(_00277_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08235_ (.I0(\as2650.stack[5][1] ),
    .I1(_02625_),
    .S(_02738_),
    .Z(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08236_ (.I(_02740_),
    .Z(_00278_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08237_ (.I0(\as2650.stack[5][2] ),
    .I1(_02627_),
    .S(_02738_),
    .Z(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08238_ (.I(_02741_),
    .Z(_00279_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08239_ (.I0(\as2650.stack[5][3] ),
    .I1(_02629_),
    .S(_02738_),
    .Z(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08240_ (.I(_02742_),
    .Z(_00280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08241_ (.I(_02737_),
    .Z(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08242_ (.I0(\as2650.stack[5][4] ),
    .I1(_02631_),
    .S(_02743_),
    .Z(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08243_ (.I(_02744_),
    .Z(_00281_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08244_ (.I0(\as2650.stack[5][5] ),
    .I1(_02634_),
    .S(_02743_),
    .Z(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08245_ (.I(_02745_),
    .Z(_00282_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08246_ (.I0(\as2650.stack[5][6] ),
    .I1(_02636_),
    .S(_02743_),
    .Z(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08247_ (.I(_02746_),
    .Z(_00283_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08248_ (.I0(\as2650.stack[5][7] ),
    .I1(_02638_),
    .S(_02743_),
    .Z(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08249_ (.I(_02747_),
    .Z(_00284_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08250_ (.I(_02737_),
    .Z(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08251_ (.I0(\as2650.stack[5][8] ),
    .I1(_02640_),
    .S(_02748_),
    .Z(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08252_ (.I(_02749_),
    .Z(_00285_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08253_ (.I0(\as2650.stack[5][9] ),
    .I1(_02643_),
    .S(_02748_),
    .Z(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08254_ (.I(_02750_),
    .Z(_00286_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08255_ (.I0(\as2650.stack[5][10] ),
    .I1(_02645_),
    .S(_02748_),
    .Z(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08256_ (.I(_02751_),
    .Z(_00287_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08257_ (.I0(\as2650.stack[5][11] ),
    .I1(_02647_),
    .S(_02748_),
    .Z(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08258_ (.I(_02752_),
    .Z(_00288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08259_ (.I(_02737_),
    .Z(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08260_ (.I0(\as2650.stack[5][12] ),
    .I1(_02649_),
    .S(_02753_),
    .Z(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08261_ (.I(_02754_),
    .Z(_00289_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08262_ (.I0(\as2650.stack[5][13] ),
    .I1(_02652_),
    .S(_02753_),
    .Z(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08263_ (.I(_02755_),
    .Z(_00290_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08264_ (.I0(\as2650.stack[5][14] ),
    .I1(_02654_),
    .S(_02753_),
    .Z(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08265_ (.I(_02756_),
    .Z(_00291_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08266_ (.I0(\as2650.stack[5][15] ),
    .I1(_02656_),
    .S(_02753_),
    .Z(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08267_ (.I(_02757_),
    .Z(_00292_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08268_ (.A1(_02247_),
    .A2(_02248_),
    .A3(_02556_),
    .A4(_02482_),
    .ZN(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08269_ (.I(_02758_),
    .Z(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08270_ (.I0(_02658_),
    .I1(\as2650.stack[10][0] ),
    .S(_02759_),
    .Z(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08271_ (.I(_02760_),
    .Z(_00293_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08272_ (.I0(_02662_),
    .I1(\as2650.stack[10][1] ),
    .S(_02759_),
    .Z(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08273_ (.I(_02761_),
    .Z(_00294_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08274_ (.I0(_02664_),
    .I1(\as2650.stack[10][2] ),
    .S(_02759_),
    .Z(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08275_ (.I(_02762_),
    .Z(_00295_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08276_ (.I0(_02666_),
    .I1(\as2650.stack[10][3] ),
    .S(_02759_),
    .Z(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08277_ (.I(_02763_),
    .Z(_00296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08278_ (.I(_02758_),
    .Z(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08279_ (.I0(_02668_),
    .I1(\as2650.stack[10][4] ),
    .S(_02764_),
    .Z(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08280_ (.I(_02765_),
    .Z(_00297_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08281_ (.I0(_02671_),
    .I1(\as2650.stack[10][5] ),
    .S(_02764_),
    .Z(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08282_ (.I(_02766_),
    .Z(_00298_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08283_ (.I0(_02673_),
    .I1(\as2650.stack[10][6] ),
    .S(_02764_),
    .Z(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08284_ (.I(_02767_),
    .Z(_00299_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08285_ (.I0(_02675_),
    .I1(\as2650.stack[10][7] ),
    .S(_02764_),
    .Z(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08286_ (.I(_02768_),
    .Z(_00300_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08287_ (.I(_02758_),
    .Z(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08288_ (.I0(_02677_),
    .I1(\as2650.stack[10][8] ),
    .S(_02769_),
    .Z(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08289_ (.I(_02770_),
    .Z(_00301_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08290_ (.I0(_02680_),
    .I1(\as2650.stack[10][9] ),
    .S(_02769_),
    .Z(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08291_ (.I(_02771_),
    .Z(_00302_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08292_ (.I0(_02682_),
    .I1(\as2650.stack[10][10] ),
    .S(_02769_),
    .Z(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08293_ (.I(_02772_),
    .Z(_00303_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08294_ (.I0(_02684_),
    .I1(\as2650.stack[10][11] ),
    .S(_02769_),
    .Z(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08295_ (.I(_02773_),
    .Z(_00304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08296_ (.I(_02758_),
    .Z(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08297_ (.I0(_02686_),
    .I1(\as2650.stack[10][12] ),
    .S(_02774_),
    .Z(_02775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08298_ (.I(_02775_),
    .Z(_00305_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08299_ (.I0(_02689_),
    .I1(\as2650.stack[10][13] ),
    .S(_02774_),
    .Z(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08300_ (.I(_02776_),
    .Z(_00306_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08301_ (.I0(_02691_),
    .I1(\as2650.stack[10][14] ),
    .S(_02774_),
    .Z(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08302_ (.I(_02777_),
    .Z(_00307_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08303_ (.I0(_02693_),
    .I1(\as2650.stack[10][15] ),
    .S(_02774_),
    .Z(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08304_ (.I(_02778_),
    .Z(_00308_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08305_ (.A1(_02246_),
    .A2(_02426_),
    .A3(_02485_),
    .A4(_02532_),
    .ZN(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08306_ (.I(_02779_),
    .Z(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08307_ (.I0(\as2650.stack[4][0] ),
    .I1(_02621_),
    .S(_02780_),
    .Z(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08308_ (.I(_02781_),
    .Z(_00309_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08309_ (.I0(\as2650.stack[4][1] ),
    .I1(_02625_),
    .S(_02780_),
    .Z(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08310_ (.I(_02782_),
    .Z(_00310_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08311_ (.I0(\as2650.stack[4][2] ),
    .I1(_02627_),
    .S(_02780_),
    .Z(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08312_ (.I(_02783_),
    .Z(_00311_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08313_ (.I0(\as2650.stack[4][3] ),
    .I1(_02629_),
    .S(_02780_),
    .Z(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08314_ (.I(_02784_),
    .Z(_00312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08315_ (.I(_02779_),
    .Z(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08316_ (.I0(\as2650.stack[4][4] ),
    .I1(_02631_),
    .S(_02785_),
    .Z(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08317_ (.I(_02786_),
    .Z(_00313_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08318_ (.I0(\as2650.stack[4][5] ),
    .I1(_02634_),
    .S(_02785_),
    .Z(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08319_ (.I(_02787_),
    .Z(_00314_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08320_ (.I0(\as2650.stack[4][6] ),
    .I1(_02636_),
    .S(_02785_),
    .Z(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08321_ (.I(_02788_),
    .Z(_00315_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08322_ (.I0(\as2650.stack[4][7] ),
    .I1(_02638_),
    .S(_02785_),
    .Z(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08323_ (.I(_02789_),
    .Z(_00316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08324_ (.I(_02779_),
    .Z(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08325_ (.I0(\as2650.stack[4][8] ),
    .I1(_02640_),
    .S(_02790_),
    .Z(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08326_ (.I(_02791_),
    .Z(_00317_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08327_ (.I0(\as2650.stack[4][9] ),
    .I1(_02643_),
    .S(_02790_),
    .Z(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08328_ (.I(_02792_),
    .Z(_00318_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08329_ (.I0(\as2650.stack[4][10] ),
    .I1(_02645_),
    .S(_02790_),
    .Z(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08330_ (.I(_02793_),
    .Z(_00319_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08331_ (.I0(\as2650.stack[4][11] ),
    .I1(_02647_),
    .S(_02790_),
    .Z(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08332_ (.I(_02794_),
    .Z(_00320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08333_ (.I(_02779_),
    .Z(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08334_ (.I0(\as2650.stack[4][12] ),
    .I1(_02649_),
    .S(_02795_),
    .Z(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08335_ (.I(_02796_),
    .Z(_00321_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08336_ (.I0(\as2650.stack[4][13] ),
    .I1(_02652_),
    .S(_02795_),
    .Z(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08337_ (.I(_02797_),
    .Z(_00322_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08338_ (.I0(\as2650.stack[4][14] ),
    .I1(_02654_),
    .S(_02795_),
    .Z(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08339_ (.I(_02798_),
    .Z(_00323_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08340_ (.I0(\as2650.stack[4][15] ),
    .I1(_02656_),
    .S(_02795_),
    .Z(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08341_ (.I(_02799_),
    .Z(_00324_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08342_ (.A1(_02405_),
    .A2(_02248_),
    .A3(_02255_),
    .A4(_02556_),
    .ZN(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08343_ (.I(_02800_),
    .Z(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08344_ (.I0(_02658_),
    .I1(\as2650.stack[15][0] ),
    .S(_02801_),
    .Z(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08345_ (.I(_02802_),
    .Z(_00325_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08346_ (.I0(_02662_),
    .I1(\as2650.stack[15][1] ),
    .S(_02801_),
    .Z(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08347_ (.I(_02803_),
    .Z(_00326_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08348_ (.I0(_02664_),
    .I1(\as2650.stack[15][2] ),
    .S(_02801_),
    .Z(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08349_ (.I(_02804_),
    .Z(_00327_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08350_ (.I0(_02666_),
    .I1(\as2650.stack[15][3] ),
    .S(_02801_),
    .Z(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08351_ (.I(_02805_),
    .Z(_00328_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08352_ (.I(_02800_),
    .Z(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08353_ (.I0(_02668_),
    .I1(\as2650.stack[15][4] ),
    .S(_02806_),
    .Z(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08354_ (.I(_02807_),
    .Z(_00329_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08355_ (.I0(_02671_),
    .I1(\as2650.stack[15][5] ),
    .S(_02806_),
    .Z(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08356_ (.I(_02808_),
    .Z(_00330_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08357_ (.I0(_02673_),
    .I1(\as2650.stack[15][6] ),
    .S(_02806_),
    .Z(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08358_ (.I(_02809_),
    .Z(_00331_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08359_ (.I0(_02675_),
    .I1(\as2650.stack[15][7] ),
    .S(_02806_),
    .Z(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08360_ (.I(_02810_),
    .Z(_00332_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08361_ (.I(_02800_),
    .Z(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08362_ (.I0(_02677_),
    .I1(\as2650.stack[15][8] ),
    .S(_02811_),
    .Z(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08363_ (.I(_02812_),
    .Z(_00333_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08364_ (.I0(_02680_),
    .I1(\as2650.stack[15][9] ),
    .S(_02811_),
    .Z(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08365_ (.I(_02813_),
    .Z(_00334_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08366_ (.I0(_02682_),
    .I1(\as2650.stack[15][10] ),
    .S(_02811_),
    .Z(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08367_ (.I(_02814_),
    .Z(_00335_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08368_ (.I0(_02684_),
    .I1(\as2650.stack[15][11] ),
    .S(_02811_),
    .Z(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08369_ (.I(_02815_),
    .Z(_00336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08370_ (.I(_02800_),
    .Z(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08371_ (.I0(_02686_),
    .I1(\as2650.stack[15][12] ),
    .S(_02816_),
    .Z(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08372_ (.I(_02817_),
    .Z(_00337_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08373_ (.I0(_02689_),
    .I1(\as2650.stack[15][13] ),
    .S(_02816_),
    .Z(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08374_ (.I(_02818_),
    .Z(_00338_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08375_ (.I0(_02691_),
    .I1(\as2650.stack[15][14] ),
    .S(_02816_),
    .Z(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08376_ (.I(_02819_),
    .Z(_00339_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08377_ (.I0(_02693_),
    .I1(\as2650.stack[15][15] ),
    .S(_02816_),
    .Z(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08378_ (.I(_02820_),
    .Z(_00340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08379_ (.I(_00803_),
    .Z(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08380_ (.I(_02821_),
    .Z(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08381_ (.I(_02822_),
    .Z(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08382_ (.I(_02823_),
    .Z(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08383_ (.I(_01476_),
    .Z(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08384_ (.I(_00785_),
    .Z(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08385_ (.I(_02826_),
    .Z(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08386_ (.I(_02827_),
    .Z(_02828_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08387_ (.I(_02828_),
    .Z(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08388_ (.A1(_02145_),
    .A2(_02210_),
    .ZN(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08389_ (.A1(_02156_),
    .A2(_02830_),
    .ZN(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08390_ (.A1(_01406_),
    .A2(_01662_),
    .ZN(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08391_ (.I(_02832_),
    .Z(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08392_ (.A1(_01503_),
    .A2(_00698_),
    .A3(_02211_),
    .A4(_02833_),
    .ZN(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08393_ (.A1(_01398_),
    .A2(_01410_),
    .Z(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08394_ (.I(_02835_),
    .ZN(_02836_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08395_ (.A1(_02834_),
    .A2(_02836_),
    .ZN(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08396_ (.A1(_01441_),
    .A2(_01469_),
    .ZN(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08397_ (.A1(_02838_),
    .A2(_02157_),
    .ZN(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08398_ (.I(_02839_),
    .Z(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08399_ (.A1(_01400_),
    .A2(_02212_),
    .A3(_02832_),
    .ZN(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08400_ (.I(_02841_),
    .Z(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08401_ (.A1(_02840_),
    .A2(_02842_),
    .ZN(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08402_ (.A1(_01503_),
    .A2(_01443_),
    .A3(_01470_),
    .A4(_01510_),
    .ZN(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08403_ (.I(_02844_),
    .Z(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08404_ (.I(_01508_),
    .Z(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08405_ (.A1(_02212_),
    .A2(_02846_),
    .A3(_01390_),
    .ZN(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08406_ (.A1(_00725_),
    .A2(_01366_),
    .A3(_01662_),
    .A4(_02847_),
    .ZN(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08407_ (.A1(_01505_),
    .A2(_02211_),
    .A3(_01510_),
    .ZN(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08408_ (.A1(_02845_),
    .A2(_02848_),
    .A3(_02849_),
    .ZN(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08409_ (.A1(_02831_),
    .A2(_02837_),
    .A3(_02843_),
    .A4(_02850_),
    .ZN(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08410_ (.A1(_02234_),
    .A2(_02851_),
    .ZN(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08411_ (.A1(_01224_),
    .A2(_01345_),
    .ZN(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08412_ (.A1(_00728_),
    .A2(_01430_),
    .A3(_02853_),
    .Z(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08413_ (.I(_00646_),
    .Z(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08414_ (.A1(_02855_),
    .A2(_01244_),
    .ZN(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08415_ (.A1(_02143_),
    .A2(_01385_),
    .A3(_02856_),
    .ZN(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08416_ (.A1(_01444_),
    .A2(_02857_),
    .Z(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08417_ (.A1(_01350_),
    .A2(_02858_),
    .ZN(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08418_ (.A1(_02152_),
    .A2(_01359_),
    .A3(_01361_),
    .A4(_01382_),
    .ZN(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08419_ (.A1(_01350_),
    .A2(_02860_),
    .ZN(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08420_ (.A1(_02854_),
    .A2(_02859_),
    .A3(_02861_),
    .ZN(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08421_ (.A1(_01345_),
    .A2(_02144_),
    .ZN(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08422_ (.A1(_00652_),
    .A2(_02833_),
    .ZN(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08423_ (.I(_00725_),
    .Z(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08424_ (.A1(_02865_),
    .A2(_00707_),
    .A3(_01399_),
    .ZN(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08425_ (.A1(_01504_),
    .A2(_02847_),
    .Z(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08426_ (.I(_02867_),
    .Z(_02868_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08427_ (.A1(_01409_),
    .A2(_01411_),
    .A3(_02866_),
    .A4(_02868_),
    .Z(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08428_ (.A1(_01430_),
    .A2(_02863_),
    .A3(_02864_),
    .A4(_02869_),
    .ZN(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08429_ (.I(_02870_),
    .Z(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08430_ (.I(_02871_),
    .Z(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08431_ (.I(_02150_),
    .Z(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08432_ (.A1(_02153_),
    .A2(_01351_),
    .A3(_02199_),
    .ZN(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08433_ (.A1(_02149_),
    .A2(_01655_),
    .ZN(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08434_ (.A1(_01665_),
    .A2(_01675_),
    .ZN(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08435_ (.A1(_02875_),
    .A2(_02876_),
    .ZN(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08436_ (.A1(_02873_),
    .A2(_02874_),
    .A3(_02877_),
    .ZN(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08437_ (.A1(_02852_),
    .A2(_02862_),
    .A3(_02872_),
    .A4(_02878_),
    .ZN(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08438_ (.A1(_02825_),
    .A2(_02829_),
    .A3(_02879_),
    .Z(_02880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08439_ (.A1(_02824_),
    .A2(_02880_),
    .ZN(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08440_ (.I(_02881_),
    .Z(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08441_ (.I(_02859_),
    .Z(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08442_ (.I(_01418_),
    .Z(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08443_ (.A1(net1),
    .A2(_02884_),
    .ZN(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08444_ (.I(_01422_),
    .Z(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08445_ (.I(_01425_),
    .Z(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08446_ (.A1(net17),
    .A2(_02886_),
    .B1(_02887_),
    .B2(net9),
    .ZN(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08447_ (.A1(_02885_),
    .A2(_02888_),
    .ZN(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08448_ (.A1(_00750_),
    .A2(_01367_),
    .B(_00751_),
    .ZN(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08449_ (.I(_02890_),
    .Z(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08450_ (.I(_02891_),
    .Z(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08451_ (.I(_02861_),
    .Z(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08452_ (.A1(_02892_),
    .A2(_02893_),
    .ZN(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08453_ (.I(_02849_),
    .Z(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08454_ (.A1(_02233_),
    .A2(_02895_),
    .ZN(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08455_ (.I(_02896_),
    .Z(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08456_ (.I(_00781_),
    .Z(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08457_ (.A1(_01458_),
    .A2(_01802_),
    .ZN(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08458_ (.A1(_01802_),
    .A2(_02898_),
    .B(_02899_),
    .ZN(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08459_ (.I(_02896_),
    .Z(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08460_ (.A1(_02233_),
    .A2(_02845_),
    .Z(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08461_ (.I(_02902_),
    .Z(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08462_ (.I(_02185_),
    .Z(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08463_ (.A1(_02232_),
    .A2(_02848_),
    .ZN(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08464_ (.I(_02905_),
    .Z(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08465_ (.A1(_02259_),
    .A2(_02837_),
    .Z(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08466_ (.I(_02907_),
    .Z(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08467_ (.I(_02905_),
    .Z(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08468_ (.A1(_02186_),
    .A2(_02909_),
    .ZN(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08469_ (.A1(_02904_),
    .A2(_02906_),
    .B(_02908_),
    .C(_02910_),
    .ZN(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08470_ (.I(_02835_),
    .Z(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08471_ (.A1(_02260_),
    .A2(_02912_),
    .ZN(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08472_ (.I(_02913_),
    .Z(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08473_ (.A1(_01325_),
    .A2(_02914_),
    .B(_02902_),
    .ZN(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08474_ (.A1(_01558_),
    .A2(_02903_),
    .B1(_02911_),
    .B2(_02915_),
    .ZN(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08475_ (.A1(_02901_),
    .A2(_02916_),
    .ZN(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08476_ (.I(_02870_),
    .Z(_02918_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08477_ (.A1(_02897_),
    .A2(_02900_),
    .B(_02917_),
    .C(_02918_),
    .ZN(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08478_ (.A1(_02890_),
    .A2(_01394_),
    .ZN(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _08479_ (.A1(_01394_),
    .A2(_01543_),
    .A3(_01549_),
    .B(_02920_),
    .ZN(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08480_ (.A1(_01323_),
    .A2(_01372_),
    .ZN(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _08481_ (.A1(_01372_),
    .A2(_01543_),
    .A3(_01549_),
    .B(_02922_),
    .ZN(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08482_ (.A1(_02921_),
    .A2(_02923_),
    .Z(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08483_ (.I(_02924_),
    .Z(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08484_ (.I(\as2650.debug_psl[3] ),
    .ZN(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08485_ (.A1(_01457_),
    .A2(_02926_),
    .ZN(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08486_ (.A1(_02206_),
    .A2(_01363_),
    .ZN(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08487_ (.A1(_02925_),
    .A2(_02927_),
    .B(_02928_),
    .ZN(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08488_ (.A1(_02925_),
    .A2(_02927_),
    .B(_02929_),
    .ZN(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08489_ (.I(_02926_),
    .Z(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08490_ (.A1(\as2650.debug_psl[0] ),
    .A2(_02931_),
    .ZN(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08491_ (.A1(_02925_),
    .A2(_02932_),
    .ZN(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08492_ (.A1(_02925_),
    .A2(_02932_),
    .Z(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08493_ (.A1(_02838_),
    .A2(_01363_),
    .ZN(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08494_ (.I(_02935_),
    .Z(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08495_ (.A1(_02933_),
    .A2(_02934_),
    .A3(_02936_),
    .ZN(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08496_ (.A1(_01357_),
    .A2(_01469_),
    .A3(_01363_),
    .ZN(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08497_ (.A1(_01403_),
    .A2(_02938_),
    .ZN(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08498_ (.I(_02939_),
    .Z(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08499_ (.A1(_02921_),
    .A2(_02923_),
    .Z(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08500_ (.A1(_02846_),
    .A2(_02941_),
    .ZN(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08501_ (.A1(_02921_),
    .A2(_02923_),
    .B(_01358_),
    .ZN(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08502_ (.A1(_01470_),
    .A2(_02941_),
    .B(_02942_),
    .C(_02943_),
    .ZN(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08503_ (.A1(_02921_),
    .A2(_02940_),
    .B(_02944_),
    .ZN(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08504_ (.A1(_02930_),
    .A2(_02937_),
    .A3(_02945_),
    .ZN(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08505_ (.I(_02946_),
    .Z(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08506_ (.I(_02870_),
    .Z(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08507_ (.A1(_02947_),
    .A2(_02948_),
    .ZN(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08508_ (.A1(_02854_),
    .A2(_02949_),
    .ZN(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08509_ (.A1(_01254_),
    .A2(_02854_),
    .B1(_02919_),
    .B2(_02950_),
    .ZN(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08510_ (.A1(_02861_),
    .A2(_02951_),
    .Z(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08511_ (.A1(_02894_),
    .A2(_02952_),
    .B(_02883_),
    .ZN(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08512_ (.A1(_02883_),
    .A2(_02889_),
    .B(_02953_),
    .ZN(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08513_ (.I(_02954_),
    .Z(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08514_ (.I(_02955_),
    .Z(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08515_ (.I(_02947_),
    .Z(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08516_ (.A1(_01409_),
    .A2(_01411_),
    .A3(_02866_),
    .A4(_02867_),
    .ZN(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08517_ (.I(_02958_),
    .Z(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08518_ (.I(_02853_),
    .Z(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _08519_ (.I(_02960_),
    .ZN(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08520_ (.A1(_01352_),
    .A2(_01563_),
    .A3(_02959_),
    .A4(_02961_),
    .ZN(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _08521_ (.A1(_02829_),
    .A2(_02962_),
    .ZN(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08522_ (.A1(_01813_),
    .A2(_02823_),
    .ZN(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08523_ (.A1(_02963_),
    .A2(_02964_),
    .ZN(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08524_ (.I(_02965_),
    .Z(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08525_ (.I(_01352_),
    .Z(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _08526_ (.A1(_02824_),
    .A2(_02880_),
    .B(_02965_),
    .C(_02967_),
    .ZN(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08527_ (.I(_02968_),
    .Z(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08528_ (.A1(_02957_),
    .A2(_02966_),
    .B1(_02969_),
    .B2(\as2650.regs[7][0] ),
    .ZN(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08529_ (.A1(_02882_),
    .A2(_02956_),
    .B(_02970_),
    .ZN(_00341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08530_ (.A1(net18),
    .A2(_01423_),
    .ZN(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08531_ (.A1(net2),
    .A2(_01419_),
    .B1(_01426_),
    .B2(net10),
    .ZN(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08532_ (.A1(_02883_),
    .A2(_02971_),
    .A3(_02972_),
    .ZN(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08533_ (.A1(_00760_),
    .A2(_01367_),
    .ZN(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08534_ (.A1(net31),
    .A2(_01416_),
    .B(_02974_),
    .ZN(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08535_ (.I(_02975_),
    .Z(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08536_ (.I(_02976_),
    .Z(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08537_ (.A1(_01356_),
    .A2(_01444_),
    .A3(_01383_),
    .ZN(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08538_ (.A1(_01431_),
    .A2(_02978_),
    .ZN(_02979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08539_ (.I(_02979_),
    .Z(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08540_ (.A1(_00728_),
    .A2(_01430_),
    .A3(_02960_),
    .ZN(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08541_ (.I(_02981_),
    .Z(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08542_ (.I(_01372_),
    .Z(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08543_ (.A1(_02975_),
    .A2(_02983_),
    .ZN(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08544_ (.A1(_01562_),
    .A2(_01566_),
    .B(_01395_),
    .ZN(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08545_ (.A1(_01564_),
    .A2(_01395_),
    .ZN(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08546_ (.A1(_01562_),
    .A2(_01566_),
    .B(_02983_),
    .ZN(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08547_ (.A1(_02984_),
    .A2(_02985_),
    .B1(_02986_),
    .B2(_02987_),
    .ZN(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08548_ (.I(_02988_),
    .Z(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08549_ (.A1(_01568_),
    .A2(_02984_),
    .A3(_02986_),
    .Z(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08550_ (.A1(_01396_),
    .A2(_01550_),
    .B(_02920_),
    .C(_02923_),
    .ZN(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08551_ (.A1(_02989_),
    .A2(_02990_),
    .B1(_02991_),
    .B2(_02934_),
    .ZN(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08552_ (.A1(_02989_),
    .A2(_02990_),
    .ZN(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08553_ (.A1(_02934_),
    .A2(_02991_),
    .ZN(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08554_ (.A1(_02993_),
    .A2(_02994_),
    .B(_02935_),
    .ZN(_02995_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08555_ (.A1(_02992_),
    .A2(_02995_),
    .ZN(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08556_ (.I(_02928_),
    .Z(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08557_ (.A1(_02924_),
    .A2(_02927_),
    .B(_02941_),
    .ZN(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08558_ (.A1(_02993_),
    .A2(_02998_),
    .ZN(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08559_ (.A1(_02984_),
    .A2(_02985_),
    .Z(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08560_ (.A1(_02939_),
    .A2(_03000_),
    .ZN(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08561_ (.A1(_01567_),
    .A2(_02984_),
    .A3(_02986_),
    .ZN(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08562_ (.A1(_01364_),
    .A2(_02989_),
    .B(_03002_),
    .C(_01442_),
    .ZN(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08563_ (.A1(_01462_),
    .A2(_02989_),
    .B(_03003_),
    .ZN(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08564_ (.A1(_02997_),
    .A2(_02999_),
    .B(_03001_),
    .C(_03004_),
    .ZN(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08565_ (.A1(_02996_),
    .A2(_03005_),
    .Z(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08566_ (.I(_03006_),
    .Z(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08567_ (.I(_02845_),
    .Z(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08568_ (.A1(_02233_),
    .A2(_03008_),
    .ZN(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08569_ (.I(_03009_),
    .Z(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08570_ (.A1(_02260_),
    .A2(_02843_),
    .ZN(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08571_ (.I(_03011_),
    .Z(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08572_ (.I(_03012_),
    .Z(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08573_ (.A1(_02189_),
    .A2(_02906_),
    .ZN(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08574_ (.A1(_02232_),
    .A2(_02848_),
    .Z(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08575_ (.I(_03015_),
    .Z(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08576_ (.A1(_02260_),
    .A2(_02837_),
    .ZN(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08577_ (.A1(_01023_),
    .A2(_03016_),
    .B(_03017_),
    .ZN(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08578_ (.A1(net182),
    .A2(_02914_),
    .B1(_03014_),
    .B2(_03018_),
    .ZN(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08579_ (.I(_03011_),
    .Z(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08580_ (.A1(_01465_),
    .A2(_01023_),
    .ZN(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08581_ (.A1(_01826_),
    .A2(_01557_),
    .ZN(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08582_ (.A1(_03020_),
    .A2(_03021_),
    .A3(_03022_),
    .ZN(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08583_ (.A1(_03013_),
    .A2(_03019_),
    .B(_03023_),
    .C(_03009_),
    .ZN(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08584_ (.A1(_01578_),
    .A2(_03010_),
    .B(_03024_),
    .C(_02901_),
    .ZN(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08585_ (.A1(_02904_),
    .A2(_02897_),
    .B(_03025_),
    .C(_02918_),
    .ZN(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08586_ (.A1(_02872_),
    .A2(_03007_),
    .B(_03026_),
    .ZN(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08587_ (.A1(_02982_),
    .A2(_03027_),
    .ZN(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08588_ (.A1(_01256_),
    .A2(_02982_),
    .B(_02980_),
    .C(_03028_),
    .ZN(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08589_ (.I(_02858_),
    .Z(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _08590_ (.A1(_01351_),
    .A2(_03030_),
    .Z(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08591_ (.I(_03031_),
    .Z(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08592_ (.A1(_02977_),
    .A2(_02980_),
    .B(_03029_),
    .C(_03032_),
    .ZN(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08593_ (.A1(_02973_),
    .A2(_03033_),
    .ZN(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08594_ (.I(_03034_),
    .Z(_03035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08595_ (.I(_02968_),
    .Z(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08596_ (.I(_03007_),
    .Z(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08597_ (.I(_02965_),
    .Z(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08598_ (.A1(\as2650.regs[7][1] ),
    .A2(_03036_),
    .B1(_03037_),
    .B2(_03038_),
    .ZN(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08599_ (.A1(_02882_),
    .A2(_03035_),
    .B(_03039_),
    .ZN(_00342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _08600_ (.A1(net3),
    .A2(_01418_),
    .B1(_02886_),
    .B2(net19),
    .C1(net11),
    .C2(_02887_),
    .ZN(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08601_ (.A1(_02883_),
    .A2(_03040_),
    .ZN(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08602_ (.I(_01369_),
    .Z(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08603_ (.A1(_01579_),
    .A2(_01052_),
    .B(_01580_),
    .ZN(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08604_ (.I(_02981_),
    .Z(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08605_ (.I(_02871_),
    .Z(_03045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08606_ (.A1(_02986_),
    .A2(_02987_),
    .ZN(_03046_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08607_ (.A1(_03000_),
    .A2(_03046_),
    .ZN(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08608_ (.I(_01394_),
    .Z(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08609_ (.I(_00715_),
    .Z(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08610_ (.A1(_03049_),
    .A2(_03048_),
    .ZN(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08611_ (.A1(_03048_),
    .A2(_01583_),
    .B(_03050_),
    .ZN(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08612_ (.I0(_02291_),
    .I1(_01583_),
    .S(_01395_),
    .Z(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08613_ (.I(_03052_),
    .Z(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08614_ (.A1(_03051_),
    .A2(_03053_),
    .Z(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08615_ (.A1(_02992_),
    .A2(_03047_),
    .B(_03054_),
    .ZN(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08616_ (.A1(_02992_),
    .A2(_03054_),
    .A3(_03047_),
    .Z(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08617_ (.A1(_02936_),
    .A2(_03055_),
    .A3(_03056_),
    .ZN(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08618_ (.I0(_01369_),
    .I1(_01583_),
    .S(_02983_),
    .Z(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08619_ (.A1(_03058_),
    .A2(_03052_),
    .Z(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08620_ (.A1(_03002_),
    .A2(_02998_),
    .B(_02988_),
    .ZN(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08621_ (.A1(_03059_),
    .A2(_03060_),
    .Z(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08622_ (.A1(_02839_),
    .A2(_03061_),
    .ZN(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08623_ (.A1(_02940_),
    .A2(_03051_),
    .ZN(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08624_ (.A1(_03058_),
    .A2(_03053_),
    .ZN(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08625_ (.A1(_01470_),
    .A2(_03064_),
    .ZN(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08626_ (.A1(_03058_),
    .A2(_03053_),
    .B(_01442_),
    .ZN(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08627_ (.A1(_02158_),
    .A2(_03064_),
    .B(_03065_),
    .C(_03066_),
    .ZN(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08628_ (.A1(_03057_),
    .A2(_03062_),
    .A3(_03063_),
    .A4(_03067_),
    .ZN(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08629_ (.I(_03068_),
    .Z(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08630_ (.I(_02896_),
    .Z(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08631_ (.I(_02902_),
    .Z(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08632_ (.A1(_01578_),
    .A2(_03021_),
    .Z(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08633_ (.I(_02913_),
    .Z(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08634_ (.A1(net193),
    .A2(_03073_),
    .B(_03011_),
    .ZN(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08635_ (.A1(_02184_),
    .A2(_02909_),
    .ZN(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08636_ (.A1(_01575_),
    .A2(_02906_),
    .B(_02908_),
    .C(_03075_),
    .ZN(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08637_ (.A1(_03020_),
    .A2(_03072_),
    .B1(_03074_),
    .B2(_03076_),
    .ZN(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08638_ (.A1(_01589_),
    .A2(_02903_),
    .ZN(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08639_ (.A1(_03071_),
    .A2(_03077_),
    .B(_03078_),
    .C(_02901_),
    .ZN(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08640_ (.A1(_01558_),
    .A2(_03070_),
    .B(_03079_),
    .C(_02948_),
    .ZN(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08641_ (.A1(_03045_),
    .A2(_03069_),
    .B(_03080_),
    .ZN(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08642_ (.A1(_03044_),
    .A2(_03081_),
    .ZN(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08643_ (.A1(_03043_),
    .A2(_02982_),
    .B(_02979_),
    .C(_03082_),
    .ZN(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08644_ (.I(_03031_),
    .Z(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08645_ (.A1(_03042_),
    .A2(_02980_),
    .B(_03083_),
    .C(_03084_),
    .ZN(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08646_ (.A1(_03041_),
    .A2(_03085_),
    .ZN(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08647_ (.I(_03086_),
    .Z(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08648_ (.I(_03087_),
    .Z(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08649_ (.I(_03069_),
    .Z(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08650_ (.A1(\as2650.regs[7][2] ),
    .A2(_03036_),
    .B1(_03089_),
    .B2(_03038_),
    .ZN(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08651_ (.A1(_02882_),
    .A2(_03088_),
    .B(_03090_),
    .ZN(_00343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _08652_ (.A1(net4),
    .A2(_02884_),
    .B1(_02886_),
    .B2(net20),
    .C1(net12),
    .C2(_02887_),
    .ZN(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08653_ (.I0(net33),
    .I1(net45),
    .S(_01416_),
    .Z(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08654_ (.I(_03092_),
    .Z(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08655_ (.I(_03093_),
    .Z(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08656_ (.A1(_03092_),
    .A2(_03048_),
    .ZN(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08657_ (.A1(_03048_),
    .A2(_01595_),
    .B(_03095_),
    .ZN(_03096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08658_ (.A1(_02940_),
    .A2(_03096_),
    .ZN(_03097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08659_ (.A1(_01342_),
    .A2(_02983_),
    .ZN(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08660_ (.A1(_01373_),
    .A2(_01595_),
    .B(_03098_),
    .ZN(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08661_ (.A1(_03096_),
    .A2(_03099_),
    .ZN(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08662_ (.A1(_03059_),
    .A2(_03060_),
    .B(_03064_),
    .ZN(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08663_ (.A1(_03100_),
    .A2(_03101_),
    .Z(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08664_ (.A1(_03100_),
    .A2(_03101_),
    .B(_02928_),
    .ZN(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08665_ (.A1(_02206_),
    .A2(_02157_),
    .ZN(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08666_ (.A1(_03096_),
    .A2(_03099_),
    .ZN(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08667_ (.I(_03105_),
    .Z(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08668_ (.A1(_01596_),
    .A2(_03095_),
    .A3(_03098_),
    .ZN(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08669_ (.A1(_03051_),
    .A2(_03053_),
    .Z(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08670_ (.A1(_03055_),
    .A2(_03106_),
    .A3(_03107_),
    .A4(_03108_),
    .Z(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08671_ (.A1(_03105_),
    .A2(_03107_),
    .B1(_03108_),
    .B2(_03055_),
    .ZN(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08672_ (.A1(_01461_),
    .A2(_03106_),
    .ZN(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08673_ (.A1(_01364_),
    .A2(_03106_),
    .ZN(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08674_ (.A1(_01358_),
    .A2(_03107_),
    .A3(_03112_),
    .ZN(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08675_ (.A1(_03104_),
    .A2(_03109_),
    .A3(_03110_),
    .B1(_03111_),
    .B2(_03113_),
    .ZN(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08676_ (.A1(_03102_),
    .A2(_03103_),
    .B(_03114_),
    .ZN(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08677_ (.A1(_03097_),
    .A2(_03115_),
    .ZN(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08678_ (.I(_03116_),
    .Z(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08679_ (.A1(_01557_),
    .A2(_01575_),
    .B(_01466_),
    .ZN(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08680_ (.A1(_01589_),
    .A2(_03118_),
    .Z(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08681_ (.A1(_02178_),
    .A2(_03015_),
    .B(_02907_),
    .ZN(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08682_ (.A1(_01073_),
    .A2(_03016_),
    .B(_03120_),
    .ZN(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08683_ (.A1(net197),
    .A2(_03073_),
    .B(_03121_),
    .ZN(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08684_ (.A1(_03020_),
    .A2(_03122_),
    .ZN(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08685_ (.A1(_03013_),
    .A2(_03119_),
    .B(_03123_),
    .C(_03071_),
    .ZN(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08686_ (.A1(_01376_),
    .A2(_01404_),
    .A3(_01509_),
    .ZN(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08687_ (.I(_03125_),
    .Z(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08688_ (.A1(_02261_),
    .A2(_03126_),
    .ZN(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08689_ (.A1(_01603_),
    .A2(_03071_),
    .B(_03124_),
    .C(_03127_),
    .ZN(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08690_ (.A1(_01576_),
    .A2(_02897_),
    .B(_02918_),
    .ZN(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08691_ (.A1(_02872_),
    .A2(_03117_),
    .B1(_03128_),
    .B2(_03129_),
    .ZN(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08692_ (.A1(_03044_),
    .A2(_03130_),
    .ZN(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08693_ (.A1(_01070_),
    .A2(_01075_),
    .ZN(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08694_ (.I(_02854_),
    .Z(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08695_ (.A1(_03132_),
    .A2(_03133_),
    .B(_02893_),
    .ZN(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08696_ (.A1(_03094_),
    .A2(_02893_),
    .B1(_03131_),
    .B2(_03134_),
    .ZN(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08697_ (.I0(_03091_),
    .I1(_03135_),
    .S(_03084_),
    .Z(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08698_ (.I(_03136_),
    .Z(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08699_ (.I(_03137_),
    .Z(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08700_ (.I(_03117_),
    .Z(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08701_ (.A1(\as2650.regs[7][3] ),
    .A2(_03036_),
    .B1(_03139_),
    .B2(_03038_),
    .ZN(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08702_ (.A1(_02882_),
    .A2(_03138_),
    .B(_03140_),
    .ZN(_00344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08703_ (.I(_02881_),
    .Z(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08704_ (.A1(net5),
    .A2(_02884_),
    .ZN(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08705_ (.A1(net21),
    .A2(_01422_),
    .B1(_01425_),
    .B2(net13),
    .ZN(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08706_ (.A1(_03142_),
    .A2(_03143_),
    .ZN(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08707_ (.I(_01086_),
    .Z(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08708_ (.I(_03145_),
    .Z(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08709_ (.I0(_01602_),
    .I1(_02180_),
    .S(_02909_),
    .Z(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08710_ (.A1(net198),
    .A2(_02914_),
    .B1(_03147_),
    .B2(_02908_),
    .C(_02902_),
    .ZN(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08711_ (.A1(_03146_),
    .A2(_02903_),
    .B(_03148_),
    .ZN(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08712_ (.A1(_01590_),
    .A2(_03127_),
    .ZN(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08713_ (.A1(_03127_),
    .A2(_03149_),
    .B(_03150_),
    .ZN(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08714_ (.A1(_00690_),
    .A2(_01416_),
    .B(_00692_),
    .ZN(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08715_ (.A1(_03152_),
    .A2(_01396_),
    .ZN(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08716_ (.A1(_01396_),
    .A2(_01608_),
    .B(_03153_),
    .ZN(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08717_ (.A1(_00638_),
    .A2(_01373_),
    .ZN(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08718_ (.A1(_01373_),
    .A2(_01608_),
    .B(_03155_),
    .ZN(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08719_ (.A1(_03154_),
    .A2(_03156_),
    .ZN(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08720_ (.I(_03157_),
    .Z(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08721_ (.A1(_03106_),
    .A2(_03102_),
    .A3(_03158_),
    .ZN(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08722_ (.A1(_03105_),
    .A2(_03102_),
    .B(_03157_),
    .ZN(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08723_ (.A1(_02997_),
    .A2(_03160_),
    .ZN(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08724_ (.A1(_03159_),
    .A2(_03161_),
    .ZN(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08725_ (.I(_03096_),
    .ZN(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08726_ (.A1(_03163_),
    .A2(_03099_),
    .Z(_03164_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08727_ (.A1(_03110_),
    .A2(_03158_),
    .A3(_03164_),
    .Z(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08728_ (.A1(_03110_),
    .A2(_03164_),
    .B(_03158_),
    .ZN(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08729_ (.A1(_02936_),
    .A2(_03165_),
    .A3(_03166_),
    .ZN(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08730_ (.I(_02939_),
    .Z(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08731_ (.I(_03154_),
    .Z(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08732_ (.A1(_03169_),
    .A2(_03156_),
    .Z(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08733_ (.A1(_02846_),
    .A2(_03170_),
    .ZN(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08734_ (.A1(_03169_),
    .A2(_03156_),
    .B(_01358_),
    .ZN(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08735_ (.A1(_01471_),
    .A2(_03170_),
    .B(_03171_),
    .C(_03172_),
    .ZN(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08736_ (.A1(_03168_),
    .A2(_03169_),
    .B(_03173_),
    .ZN(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08737_ (.A1(_03162_),
    .A2(_03167_),
    .A3(_03174_),
    .ZN(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08738_ (.I(_03175_),
    .Z(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08739_ (.A1(_02871_),
    .A2(_03176_),
    .ZN(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08740_ (.A1(_02918_),
    .A2(_03151_),
    .B(_03177_),
    .ZN(_03178_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08741_ (.I0(_01604_),
    .I1(_03178_),
    .S(_02981_),
    .Z(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08742_ (.I(_00664_),
    .Z(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08743_ (.A1(net34),
    .A2(_03180_),
    .B(_00719_),
    .ZN(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08744_ (.I(_03181_),
    .Z(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08745_ (.A1(_03182_),
    .A2(_02861_),
    .ZN(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08746_ (.A1(_02893_),
    .A2(_03179_),
    .B(_03183_),
    .ZN(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08747_ (.A1(_03084_),
    .A2(_03184_),
    .ZN(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08748_ (.A1(_03084_),
    .A2(_03144_),
    .B(_03185_),
    .ZN(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08749_ (.I(_03186_),
    .Z(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08750_ (.I(_03187_),
    .Z(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08751_ (.I(_03176_),
    .Z(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08752_ (.A1(\as2650.regs[7][4] ),
    .A2(_03036_),
    .B1(_03189_),
    .B2(_03038_),
    .ZN(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08753_ (.A1(_03141_),
    .A2(_03188_),
    .B(_03190_),
    .ZN(_00345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08754_ (.A1(net6),
    .A2(_01419_),
    .ZN(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08755_ (.A1(net22),
    .A2(_01423_),
    .B1(_01426_),
    .B2(net14),
    .ZN(_03192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08756_ (.A1(_03191_),
    .A2(_03192_),
    .ZN(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08757_ (.A1(_00695_),
    .A2(_01417_),
    .ZN(_03194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08758_ (.A1(net26),
    .A2(_01417_),
    .B(_03194_),
    .ZN(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08759_ (.I(_03195_),
    .Z(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08760_ (.I(_02979_),
    .Z(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08761_ (.I0(_03195_),
    .I1(_01624_),
    .S(_01374_),
    .Z(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08762_ (.I0(_01622_),
    .I1(_01624_),
    .S(_01397_),
    .Z(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08763_ (.A1(_03198_),
    .A2(_03199_),
    .Z(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08764_ (.A1(_03198_),
    .A2(_03199_),
    .ZN(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08765_ (.A1(_03200_),
    .A2(_03201_),
    .ZN(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08766_ (.I(_03169_),
    .ZN(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08767_ (.A1(_03203_),
    .A2(_03156_),
    .ZN(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08768_ (.A1(_03166_),
    .A2(_03202_),
    .A3(_03204_),
    .ZN(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08769_ (.A1(_03166_),
    .A2(_03204_),
    .B(_03202_),
    .ZN(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08770_ (.A1(_03104_),
    .A2(_03206_),
    .ZN(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08771_ (.A1(_03205_),
    .A2(_03207_),
    .ZN(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08772_ (.A1(_03170_),
    .A2(_03160_),
    .ZN(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08773_ (.A1(_03202_),
    .A2(_03209_),
    .ZN(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08774_ (.A1(_01471_),
    .A2(_03201_),
    .ZN(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08775_ (.A1(_02158_),
    .A2(_03201_),
    .ZN(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08776_ (.A1(_01443_),
    .A2(_03200_),
    .A3(_03212_),
    .ZN(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08777_ (.A1(_02840_),
    .A2(_03210_),
    .B1(_03211_),
    .B2(_03213_),
    .C(_03168_),
    .ZN(_03214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08778_ (.A1(_03168_),
    .A2(_03198_),
    .B1(_03208_),
    .B2(_03214_),
    .ZN(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08779_ (.I(_03215_),
    .Z(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08780_ (.I(_01633_),
    .Z(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08781_ (.I(_03217_),
    .Z(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08782_ (.I0(_03145_),
    .I1(_02175_),
    .S(_02905_),
    .Z(_03219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08783_ (.A1(net199),
    .A2(_03073_),
    .B1(_03219_),
    .B2(_02908_),
    .ZN(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08784_ (.A1(_02225_),
    .A2(_03145_),
    .Z(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08785_ (.A1(_03012_),
    .A2(_03221_),
    .ZN(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08786_ (.A1(_03012_),
    .A2(_03220_),
    .B(_03222_),
    .C(_03009_),
    .ZN(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08787_ (.A1(_03218_),
    .A2(_03010_),
    .B(_03223_),
    .C(_02901_),
    .ZN(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08788_ (.A1(_01603_),
    .A2(_03070_),
    .B(_03224_),
    .C(_02948_),
    .ZN(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08789_ (.A1(_03045_),
    .A2(_03216_),
    .B(_03225_),
    .ZN(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08790_ (.A1(_03044_),
    .A2(_03226_),
    .ZN(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08791_ (.A1(_01620_),
    .A2(_03133_),
    .ZN(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08792_ (.A1(_03197_),
    .A2(_03227_),
    .A3(_03228_),
    .ZN(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08793_ (.A1(_03196_),
    .A2(_02980_),
    .B(_03229_),
    .C(_03031_),
    .ZN(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08794_ (.A1(_03032_),
    .A2(_03193_),
    .B(_03230_),
    .ZN(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08795_ (.I(_03231_),
    .Z(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08796_ (.I(_03232_),
    .Z(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08797_ (.I(_03216_),
    .Z(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08798_ (.A1(\as2650.regs[7][5] ),
    .A2(_02969_),
    .B1(_03234_),
    .B2(_02966_),
    .ZN(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08799_ (.A1(_03141_),
    .A2(_03233_),
    .B(_03235_),
    .ZN(_00346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08800_ (.A1(net7),
    .A2(_02884_),
    .ZN(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08801_ (.A1(net23),
    .A2(_02886_),
    .B1(_02887_),
    .B2(net15),
    .ZN(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08802_ (.A1(_03236_),
    .A2(_03237_),
    .ZN(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08803_ (.A1(net27),
    .A2(_03180_),
    .B(_00704_),
    .ZN(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08804_ (.I(_03239_),
    .Z(_03240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _08805_ (.I(_03240_),
    .Z(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08806_ (.I(_02940_),
    .Z(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08807_ (.A1(_00680_),
    .A2(_01417_),
    .B(_00685_),
    .ZN(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08808_ (.A1(_01397_),
    .A2(_01637_),
    .ZN(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08809_ (.A1(_03243_),
    .A2(_01397_),
    .B(_03244_),
    .ZN(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08810_ (.I(_03245_),
    .Z(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08811_ (.A1(_01374_),
    .A2(_01637_),
    .ZN(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08812_ (.A1(_00623_),
    .A2(_01375_),
    .B(_03247_),
    .ZN(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08813_ (.A1(_03245_),
    .A2(_03248_),
    .ZN(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08814_ (.A1(_03245_),
    .A2(_03248_),
    .Z(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08815_ (.A1(_03249_),
    .A2(_03250_),
    .ZN(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08816_ (.I(_03198_),
    .ZN(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08817_ (.A1(_03252_),
    .A2(_03199_),
    .ZN(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08818_ (.A1(_03206_),
    .A2(_03251_),
    .A3(_03253_),
    .ZN(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08819_ (.I(_02936_),
    .Z(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08820_ (.A1(_03206_),
    .A2(_03253_),
    .B(_03251_),
    .ZN(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08821_ (.A1(_03255_),
    .A2(_03256_),
    .ZN(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08822_ (.A1(_03254_),
    .A2(_03257_),
    .ZN(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08823_ (.A1(_03170_),
    .A2(_03160_),
    .A3(_03201_),
    .ZN(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08824_ (.A1(_03200_),
    .A2(_03259_),
    .ZN(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08825_ (.A1(_03251_),
    .A2(_03260_),
    .Z(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08826_ (.A1(_02997_),
    .A2(_03261_),
    .ZN(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08827_ (.A1(_01471_),
    .A2(_03250_),
    .B1(_03251_),
    .B2(_01365_),
    .ZN(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08828_ (.A1(_01359_),
    .A2(_03263_),
    .ZN(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08829_ (.A1(_02211_),
    .A2(_02938_),
    .A3(_03264_),
    .ZN(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08830_ (.A1(_03258_),
    .A2(_03262_),
    .A3(_03265_),
    .ZN(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08831_ (.A1(_03242_),
    .A2(_03246_),
    .B(_03266_),
    .ZN(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08832_ (.A1(_03045_),
    .A2(_03267_),
    .Z(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08833_ (.I(_02898_),
    .Z(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08834_ (.A1(_03218_),
    .A2(_03016_),
    .ZN(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08835_ (.A1(_02173_),
    .A2(_02906_),
    .B(_03017_),
    .ZN(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08836_ (.A1(net200),
    .A2(_02914_),
    .B1(_03270_),
    .B2(_03271_),
    .ZN(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08837_ (.A1(_02225_),
    .A2(_03145_),
    .ZN(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08838_ (.A1(_03218_),
    .A2(_03273_),
    .Z(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08839_ (.A1(_03020_),
    .A2(_03274_),
    .ZN(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08840_ (.A1(_03013_),
    .A2(_03272_),
    .B(_03275_),
    .C(_03010_),
    .ZN(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08841_ (.A1(_03269_),
    .A2(_03010_),
    .B(_03276_),
    .C(_03070_),
    .ZN(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08842_ (.A1(_03146_),
    .A2(_02897_),
    .B(_03277_),
    .C(_02872_),
    .ZN(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08843_ (.A1(_03268_),
    .A2(_03278_),
    .B(_03133_),
    .ZN(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08844_ (.A1(_00988_),
    .A2(_03133_),
    .ZN(_03280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08845_ (.A1(_03197_),
    .A2(_03280_),
    .ZN(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _08846_ (.A1(_03241_),
    .A2(_03197_),
    .B1(_03279_),
    .B2(_03281_),
    .C(_03031_),
    .ZN(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08847_ (.A1(_03032_),
    .A2(_03238_),
    .B(_03282_),
    .ZN(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08848_ (.I(_03283_),
    .Z(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08849_ (.I(_03284_),
    .Z(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08850_ (.I(_03267_),
    .Z(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08851_ (.A1(\as2650.regs[7][6] ),
    .A2(_02969_),
    .B1(_03286_),
    .B2(_02966_),
    .ZN(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08852_ (.A1(_03141_),
    .A2(_03285_),
    .B(_03287_),
    .ZN(_00347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08853_ (.A1(net8),
    .A2(_01419_),
    .ZN(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08854_ (.A1(net24),
    .A2(_01423_),
    .B1(_01426_),
    .B2(net16),
    .ZN(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08855_ (.A1(_03288_),
    .A2(_03289_),
    .ZN(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08856_ (.I(_01669_),
    .Z(_03291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08857_ (.A1(_03291_),
    .A2(_02860_),
    .B(_03030_),
    .ZN(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08858_ (.A1(_01432_),
    .A2(_03292_),
    .ZN(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08859_ (.I0(_01668_),
    .I1(_01646_),
    .S(_01374_),
    .Z(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08860_ (.I0(_01644_),
    .I1(_01646_),
    .S(_01398_),
    .Z(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08861_ (.A1(_03294_),
    .A2(_03295_),
    .Z(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08862_ (.A1(_03294_),
    .A2(_03295_),
    .ZN(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08863_ (.A1(_03296_),
    .A2(_03297_),
    .ZN(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08864_ (.I(_03248_),
    .ZN(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08865_ (.A1(_03246_),
    .A2(_03299_),
    .ZN(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08866_ (.A1(_03256_),
    .A2(_03298_),
    .A3(_03300_),
    .Z(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08867_ (.A1(_03256_),
    .A2(_03300_),
    .B(_03298_),
    .ZN(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08868_ (.A1(_03104_),
    .A2(_03301_),
    .A3(_03302_),
    .Z(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08869_ (.A1(_03246_),
    .A2(_03248_),
    .Z(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _08870_ (.A1(_03200_),
    .A2(_03304_),
    .A3(_03259_),
    .B(_03250_),
    .ZN(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08871_ (.A1(_03298_),
    .A2(_03305_),
    .Z(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08872_ (.A1(_01462_),
    .A2(_03297_),
    .B1(_03298_),
    .B2(_02158_),
    .ZN(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08873_ (.A1(_01444_),
    .A2(_03307_),
    .ZN(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08874_ (.A1(_02840_),
    .A2(_03306_),
    .B(_03308_),
    .C(_03168_),
    .ZN(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08875_ (.A1(_03242_),
    .A2(_03294_),
    .B1(_03303_),
    .B2(_03309_),
    .ZN(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08876_ (.I(_03310_),
    .Z(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08877_ (.A1(_01802_),
    .A2(_02187_),
    .B(_02899_),
    .ZN(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08878_ (.A1(_03217_),
    .A2(_01616_),
    .B(_02225_),
    .ZN(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08879_ (.A1(_02898_),
    .A2(_03313_),
    .Z(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08880_ (.A1(_03269_),
    .A2(_03016_),
    .ZN(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08881_ (.A1(_02165_),
    .A2(_02909_),
    .B(_03017_),
    .ZN(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08882_ (.A1(_00619_),
    .A2(_03073_),
    .B1(_03315_),
    .B2(_03316_),
    .ZN(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08883_ (.A1(_03012_),
    .A2(_03317_),
    .ZN(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08884_ (.A1(_03013_),
    .A2(_03314_),
    .B(_03318_),
    .C(_02903_),
    .ZN(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08885_ (.A1(_03071_),
    .A2(_03312_),
    .B(_03319_),
    .C(_03127_),
    .ZN(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08886_ (.A1(_01630_),
    .A2(_03070_),
    .B(_02948_),
    .ZN(_03321_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08887_ (.A1(_03045_),
    .A2(_03311_),
    .B1(_03320_),
    .B2(_03321_),
    .ZN(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08888_ (.A1(_03044_),
    .A2(_03322_),
    .ZN(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08889_ (.A1(_01642_),
    .A2(_02982_),
    .B(_03197_),
    .C(_03323_),
    .ZN(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08890_ (.A1(_03293_),
    .A2(_03324_),
    .ZN(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08891_ (.A1(_03032_),
    .A2(_03290_),
    .B(_03325_),
    .ZN(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08892_ (.I(_03326_),
    .Z(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08893_ (.I(_03327_),
    .Z(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08894_ (.I(_03311_),
    .Z(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08895_ (.I(_03329_),
    .Z(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08896_ (.A1(\as2650.regs[7][7] ),
    .A2(_02969_),
    .B1(_03330_),
    .B2(_02966_),
    .ZN(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08897_ (.A1(_03141_),
    .A2(_03328_),
    .B(_03331_),
    .ZN(_00348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _08898_ (.A1(_02486_),
    .A2(_02599_),
    .ZN(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08899_ (.I(_03332_),
    .Z(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08900_ (.I0(_02555_),
    .I1(\as2650.stack[1][0] ),
    .S(_03333_),
    .Z(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08901_ (.I(_03334_),
    .Z(_00349_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08902_ (.I0(_02560_),
    .I1(\as2650.stack[1][1] ),
    .S(_03333_),
    .Z(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08903_ (.I(_03335_),
    .Z(_00350_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08904_ (.I0(_02562_),
    .I1(\as2650.stack[1][2] ),
    .S(_03333_),
    .Z(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08905_ (.I(_03336_),
    .Z(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08906_ (.I0(_02564_),
    .I1(\as2650.stack[1][3] ),
    .S(_03333_),
    .Z(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08907_ (.I(_03337_),
    .Z(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08908_ (.I(_03332_),
    .Z(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08909_ (.I0(_02566_),
    .I1(\as2650.stack[1][4] ),
    .S(_03338_),
    .Z(_03339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08910_ (.I(_03339_),
    .Z(_00353_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08911_ (.I0(_02569_),
    .I1(\as2650.stack[1][5] ),
    .S(_03338_),
    .Z(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08912_ (.I(_03340_),
    .Z(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08913_ (.I0(_02571_),
    .I1(\as2650.stack[1][6] ),
    .S(_03338_),
    .Z(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08914_ (.I(_03341_),
    .Z(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08915_ (.I0(_02573_),
    .I1(\as2650.stack[1][7] ),
    .S(_03338_),
    .Z(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08916_ (.I(_03342_),
    .Z(_00356_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08917_ (.I(_03332_),
    .Z(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08918_ (.I0(_02575_),
    .I1(\as2650.stack[1][8] ),
    .S(_03343_),
    .Z(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08919_ (.I(_03344_),
    .Z(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08920_ (.I0(_02578_),
    .I1(\as2650.stack[1][9] ),
    .S(_03343_),
    .Z(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08921_ (.I(_03345_),
    .Z(_00358_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08922_ (.I0(_02580_),
    .I1(\as2650.stack[1][10] ),
    .S(_03343_),
    .Z(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08923_ (.I(_03346_),
    .Z(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08924_ (.I0(_02582_),
    .I1(\as2650.stack[1][11] ),
    .S(_03343_),
    .Z(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08925_ (.I(_03347_),
    .Z(_00360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08926_ (.I(_03332_),
    .Z(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08927_ (.I0(_02584_),
    .I1(\as2650.stack[1][12] ),
    .S(_03348_),
    .Z(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08928_ (.I(_03349_),
    .Z(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08929_ (.I0(_02587_),
    .I1(\as2650.stack[1][13] ),
    .S(_03348_),
    .Z(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08930_ (.I(_03350_),
    .Z(_00362_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08931_ (.I0(_02589_),
    .I1(\as2650.stack[1][14] ),
    .S(_03348_),
    .Z(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08932_ (.I(_03351_),
    .Z(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08933_ (.I0(_02591_),
    .I1(\as2650.stack[1][15] ),
    .S(_03348_),
    .Z(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08934_ (.I(_03352_),
    .Z(_00364_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08935_ (.I(_01538_),
    .Z(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08936_ (.A1(\as2650.last_addr[0] ),
    .A2(_03353_),
    .ZN(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08937_ (.A1(_01555_),
    .A2(_03354_),
    .B(_01685_),
    .ZN(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08938_ (.A1(_01279_),
    .A2(net205),
    .ZN(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08939_ (.A1(\as2650.last_addr[1] ),
    .A2(_01539_),
    .ZN(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08940_ (.A1(_01435_),
    .A2(_03355_),
    .A3(_03356_),
    .ZN(_00366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08941_ (.I(_01684_),
    .Z(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08942_ (.A1(\as2650.last_addr[2] ),
    .A2(_01577_),
    .B(_01586_),
    .ZN(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08943_ (.A1(_03357_),
    .A2(_03358_),
    .ZN(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08944_ (.A1(_01287_),
    .A2(net205),
    .ZN(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08945_ (.A1(\as2650.last_addr[3] ),
    .A2(_03353_),
    .ZN(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08946_ (.A1(_01435_),
    .A2(_03359_),
    .A3(_03360_),
    .ZN(_00368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08947_ (.A1(_01295_),
    .A2(_01571_),
    .ZN(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08948_ (.A1(\as2650.last_addr[4] ),
    .A2(_01560_),
    .ZN(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08949_ (.A1(_03361_),
    .A2(_03362_),
    .B(_01685_),
    .ZN(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08950_ (.A1(\as2650.last_addr[5] ),
    .A2(_03353_),
    .ZN(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08951_ (.A1(_01435_),
    .A2(_01629_),
    .A3(_03363_),
    .ZN(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08952_ (.A1(_01308_),
    .A2(_01571_),
    .ZN(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08953_ (.A1(\as2650.last_addr[6] ),
    .A2(_01560_),
    .ZN(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08954_ (.A1(_03364_),
    .A2(_03365_),
    .B(_01685_),
    .ZN(_00371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08955_ (.I(_01449_),
    .Z(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08956_ (.A1(\as2650.last_addr[7] ),
    .A2(_03353_),
    .ZN(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08957_ (.A1(_03366_),
    .A2(_01651_),
    .A3(_03367_),
    .ZN(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08958_ (.I(_01529_),
    .ZN(_00374_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08959_ (.I(\as2650.indirect_target[0] ),
    .ZN(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08960_ (.I(_01348_),
    .Z(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08961_ (.I(_03369_),
    .Z(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08962_ (.I(_01684_),
    .Z(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08963_ (.A1(_01356_),
    .A2(_01385_),
    .A3(_01243_),
    .ZN(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08964_ (.I(_01657_),
    .Z(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08965_ (.I(_01674_),
    .Z(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08966_ (.A1(_03372_),
    .A2(_03373_),
    .A3(_03374_),
    .ZN(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08967_ (.I(_03375_),
    .Z(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08968_ (.I(_02207_),
    .Z(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08969_ (.A1(_03373_),
    .A2(_03374_),
    .ZN(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08970_ (.A1(_00717_),
    .A2(_03378_),
    .ZN(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08971_ (.I(_03379_),
    .ZN(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08972_ (.A1(_02207_),
    .A2(_03380_),
    .B(_01677_),
    .ZN(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08973_ (.I(_01349_),
    .Z(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _08974_ (.A1(_01343_),
    .A2(_03382_),
    .A3(_02144_),
    .B(\as2650.instruction_args_latch[8] ),
    .ZN(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08975_ (.A1(_02891_),
    .A2(_01653_),
    .A3(_01428_),
    .A4(_01386_),
    .ZN(_03384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08976_ (.A1(_03383_),
    .A2(_03384_),
    .ZN(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08977_ (.A1(_02281_),
    .A2(_03385_),
    .Z(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08978_ (.A1(_02892_),
    .A2(_03377_),
    .A3(_03379_),
    .B1(_03381_),
    .B2(_03386_),
    .ZN(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _08979_ (.A1(_02873_),
    .A2(_02876_),
    .Z(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08980_ (.I(_03388_),
    .Z(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08981_ (.A1(_01667_),
    .A2(_03387_),
    .B1(_03389_),
    .B2(_03368_),
    .ZN(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08982_ (.A1(_03372_),
    .A2(_01346_),
    .ZN(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08983_ (.I(_03391_),
    .Z(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08984_ (.I(_03378_),
    .Z(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08985_ (.A1(_03392_),
    .A2(_03393_),
    .ZN(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08986_ (.A1(_00957_),
    .A2(_01652_),
    .A3(_01428_),
    .ZN(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08987_ (.I(_03395_),
    .Z(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08988_ (.I(_03396_),
    .Z(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08989_ (.I(_03397_),
    .Z(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08990_ (.A1(_03372_),
    .A2(_02890_),
    .A3(_01343_),
    .A4(_03382_),
    .ZN(_03399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08991_ (.A1(_01008_),
    .A2(_03398_),
    .B(_03399_),
    .ZN(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08992_ (.A1(_03376_),
    .A2(_03390_),
    .B1(_03394_),
    .B2(_03400_),
    .ZN(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08993_ (.A1(_03368_),
    .A2(_03370_),
    .B(_03371_),
    .C(_03401_),
    .ZN(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08994_ (.I(\as2650.indirect_target[1] ),
    .ZN(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08995_ (.A1(_02212_),
    .A2(_03374_),
    .A3(_01675_),
    .ZN(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08996_ (.A1(_03383_),
    .A2(_03384_),
    .B(_02222_),
    .ZN(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _08997_ (.A1(_01344_),
    .A2(_03382_),
    .A3(_02144_),
    .B(\as2650.instruction_args_latch[9] ),
    .ZN(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08998_ (.A1(_00760_),
    .A2(net123),
    .B(_00761_),
    .ZN(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08999_ (.A1(_03406_),
    .A2(_01653_),
    .A3(_01429_),
    .A4(_01387_),
    .ZN(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09000_ (.A1(_03405_),
    .A2(_03407_),
    .ZN(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _09001_ (.I(_03408_),
    .ZN(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09002_ (.A1(_02282_),
    .A2(_03404_),
    .A3(_03409_),
    .Z(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09003_ (.I(_02206_),
    .Z(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09004_ (.I(_01507_),
    .Z(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09005_ (.A1(_03411_),
    .A2(_00722_),
    .A3(_03412_),
    .A4(_01659_),
    .Z(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09006_ (.I(_03413_),
    .Z(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09007_ (.A1(_03413_),
    .A2(_03410_),
    .ZN(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09008_ (.A1(_02976_),
    .A2(_03414_),
    .B(_03415_),
    .ZN(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09009_ (.I(_03379_),
    .Z(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09010_ (.A1(_03403_),
    .A2(_03410_),
    .B1(_03416_),
    .B2(_03417_),
    .ZN(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09011_ (.A1(_03402_),
    .A2(_03389_),
    .B1(_03418_),
    .B2(_01667_),
    .ZN(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _09012_ (.A1(_03372_),
    .A2(_01344_),
    .A3(_03382_),
    .B(\as2650.instruction_args_latch[1] ),
    .ZN(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _09013_ (.A1(_02149_),
    .A2(_03406_),
    .A3(_01654_),
    .A4(_01429_),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09014_ (.A1(_03420_),
    .A2(_03421_),
    .ZN(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09015_ (.I(_03394_),
    .Z(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09016_ (.A1(_03376_),
    .A2(_03419_),
    .B1(_03422_),
    .B2(_03423_),
    .ZN(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09017_ (.A1(_03402_),
    .A2(_03370_),
    .B(_03371_),
    .C(_03424_),
    .ZN(_00377_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09018_ (.I(\as2650.indirect_target[2] ),
    .ZN(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09019_ (.I(_03388_),
    .Z(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09020_ (.I0(_03049_),
    .I1(\as2650.instruction_args_latch[10] ),
    .S(_01670_),
    .Z(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09021_ (.I(_03427_),
    .Z(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09022_ (.A1(_02282_),
    .A2(_03405_),
    .A3(_03407_),
    .ZN(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09023_ (.A1(_03405_),
    .A2(_03407_),
    .B(_02282_),
    .ZN(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09024_ (.A1(_03404_),
    .A2(_03429_),
    .B(_03430_),
    .ZN(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09025_ (.A1(_02298_),
    .A2(_03428_),
    .A3(_03431_),
    .Z(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09026_ (.I(_03049_),
    .Z(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09027_ (.I0(_03433_),
    .I1(_03432_),
    .S(_02207_),
    .Z(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09028_ (.A1(_03403_),
    .A2(_03432_),
    .B1(_03434_),
    .B2(_03417_),
    .ZN(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09029_ (.A1(_03425_),
    .A2(_03426_),
    .B1(_03435_),
    .B2(_01667_),
    .ZN(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09030_ (.I0(_03049_),
    .I1(\as2650.instruction_args_latch[2] ),
    .S(_03395_),
    .Z(_03437_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09031_ (.A1(_03376_),
    .A2(_03436_),
    .B1(_03437_),
    .B2(_03423_),
    .ZN(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09032_ (.A1(_03425_),
    .A2(_03370_),
    .B(_03371_),
    .C(_03438_),
    .ZN(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09033_ (.I(\as2650.indirect_target[3] ),
    .ZN(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09034_ (.I(_01683_),
    .Z(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09035_ (.I(_03440_),
    .Z(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09036_ (.I(_01670_),
    .Z(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _09037_ (.I(\as2650.instruction_args_latch[11] ),
    .ZN(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09038_ (.A1(_03443_),
    .A2(_03442_),
    .ZN(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09039_ (.A1(_03092_),
    .A2(_03442_),
    .B(_03444_),
    .ZN(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09040_ (.A1(_02295_),
    .A2(_02297_),
    .ZN(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09041_ (.A1(_03446_),
    .A2(_03427_),
    .ZN(_03447_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09042_ (.I(_03446_),
    .Z(_03448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09043_ (.A1(_03448_),
    .A2(_03427_),
    .ZN(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09044_ (.A1(_03447_),
    .A2(_03431_),
    .B(_03449_),
    .ZN(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09045_ (.A1(_02310_),
    .A2(_03445_),
    .A3(_03450_),
    .Z(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09046_ (.A1(net33),
    .A2(_03180_),
    .B(_00710_),
    .ZN(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09047_ (.I(_03452_),
    .Z(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09048_ (.I(_03414_),
    .Z(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09049_ (.I(_03413_),
    .Z(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09050_ (.A1(_03455_),
    .A2(_03451_),
    .ZN(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09051_ (.A1(_03453_),
    .A2(_03454_),
    .B(_03456_),
    .ZN(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09052_ (.A1(_03403_),
    .A2(_03451_),
    .B1(_03457_),
    .B2(_03417_),
    .ZN(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09053_ (.I(_01666_),
    .Z(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09054_ (.A1(_03439_),
    .A2(_03426_),
    .B1(_03458_),
    .B2(_03459_),
    .ZN(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09055_ (.A1(\as2650.instruction_args_latch[3] ),
    .A2(_03395_),
    .ZN(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09056_ (.A1(_03452_),
    .A2(_03395_),
    .B(_03461_),
    .ZN(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09057_ (.I(_03394_),
    .Z(_03463_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09058_ (.A1(_03376_),
    .A2(_03460_),
    .B1(_03462_),
    .B2(_03463_),
    .ZN(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09059_ (.A1(_03439_),
    .A2(_03370_),
    .B(_03441_),
    .C(_03464_),
    .ZN(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09060_ (.I(\as2650.indirect_target[4] ),
    .ZN(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09061_ (.I(_01347_),
    .Z(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09062_ (.I(_03466_),
    .Z(_03467_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09063_ (.I(_03375_),
    .Z(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09064_ (.I(_03152_),
    .Z(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09065_ (.I(_03469_),
    .Z(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09066_ (.I(_03381_),
    .Z(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09067_ (.A1(\as2650.instruction_args_latch[12] ),
    .A2(_01671_),
    .ZN(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09068_ (.A1(_03181_),
    .A2(_03442_),
    .B(_03472_),
    .ZN(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09069_ (.A1(_02324_),
    .A2(_03473_),
    .Z(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09070_ (.A1(_02310_),
    .A2(_03445_),
    .ZN(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09071_ (.A1(_02310_),
    .A2(_03445_),
    .ZN(_03476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09072_ (.A1(_03475_),
    .A2(_03450_),
    .B(_03476_),
    .ZN(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09073_ (.A1(_03474_),
    .A2(_03477_),
    .Z(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09074_ (.A1(_03470_),
    .A2(_03377_),
    .A3(_03379_),
    .B1(_03471_),
    .B2(_03478_),
    .ZN(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09075_ (.A1(_03465_),
    .A2(_03426_),
    .B1(_03479_),
    .B2(_03459_),
    .ZN(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09076_ (.A1(\as2650.instruction_args_latch[4] ),
    .A2(_03396_),
    .ZN(_03481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09077_ (.A1(_03181_),
    .A2(_03397_),
    .B(_03481_),
    .ZN(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09078_ (.A1(_03468_),
    .A2(_03480_),
    .B1(_03482_),
    .B2(_03463_),
    .ZN(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09079_ (.A1(_03465_),
    .A2(_03467_),
    .B(_03441_),
    .C(_03483_),
    .ZN(_00380_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09080_ (.I(\as2650.indirect_target[5] ),
    .ZN(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09081_ (.A1(_02334_),
    .A2(_02337_),
    .Z(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09082_ (.I(_03442_),
    .Z(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09083_ (.A1(_00723_),
    .A2(_03486_),
    .ZN(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09084_ (.A1(_03195_),
    .A2(_03486_),
    .B(_03487_),
    .ZN(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09085_ (.A1(_02321_),
    .A2(_02323_),
    .Z(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09086_ (.I(_03473_),
    .Z(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09087_ (.A1(_03489_),
    .A2(_03490_),
    .ZN(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09088_ (.A1(_03474_),
    .A2(_03477_),
    .B(_03491_),
    .ZN(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09089_ (.A1(_03485_),
    .A2(_03488_),
    .A3(_03492_),
    .Z(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09090_ (.A1(_03455_),
    .A2(_03493_),
    .ZN(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09091_ (.A1(_03196_),
    .A2(_03454_),
    .B(_03494_),
    .ZN(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _09092_ (.A1(_03403_),
    .A2(_03493_),
    .B1(_03495_),
    .B2(_03417_),
    .ZN(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09093_ (.A1(_03484_),
    .A2(_03426_),
    .B1(_03496_),
    .B2(_03459_),
    .ZN(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09094_ (.A1(\as2650.instruction_args_latch[5] ),
    .A2(_03396_),
    .ZN(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09095_ (.A1(_03195_),
    .A2(_03397_),
    .B(_03498_),
    .ZN(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09096_ (.A1(_03468_),
    .A2(_03497_),
    .B1(_03499_),
    .B2(_03463_),
    .ZN(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09097_ (.A1(_03484_),
    .A2(_03467_),
    .B(_03441_),
    .C(_03500_),
    .ZN(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09098_ (.I(\as2650.indirect_target[6] ),
    .ZN(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09099_ (.I(_03388_),
    .Z(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09100_ (.A1(\as2650.instruction_args_latch[14] ),
    .A2(_01671_),
    .ZN(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09101_ (.A1(_03239_),
    .A2(_01671_),
    .B(_03503_),
    .ZN(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09102_ (.A1(_02353_),
    .A2(_03504_),
    .ZN(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _09103_ (.A1(_03485_),
    .A2(_03488_),
    .Z(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _09104_ (.A1(_03485_),
    .A2(_03488_),
    .Z(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09105_ (.A1(_03506_),
    .A2(_03492_),
    .B(_03507_),
    .ZN(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09106_ (.A1(_03505_),
    .A2(_03508_),
    .Z(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09107_ (.A1(_03241_),
    .A2(_03454_),
    .A3(_03380_),
    .ZN(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09108_ (.A1(_03471_),
    .A2(_03509_),
    .B(_03510_),
    .ZN(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09109_ (.A1(_03501_),
    .A2(_03502_),
    .B1(_03511_),
    .B2(_03459_),
    .ZN(_03512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09110_ (.A1(\as2650.instruction_args_latch[6] ),
    .A2(_03398_),
    .ZN(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09111_ (.A1(_03240_),
    .A2(_03398_),
    .B(_03513_),
    .ZN(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09112_ (.A1(_03468_),
    .A2(_03512_),
    .B1(_03514_),
    .B2(_03463_),
    .ZN(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09113_ (.A1(_03501_),
    .A2(_03467_),
    .B(_03441_),
    .C(_03515_),
    .ZN(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09114_ (.I(\as2650.indirect_target[7] ),
    .ZN(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09115_ (.I(_01354_),
    .Z(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09116_ (.I(_03504_),
    .Z(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09117_ (.I(_03518_),
    .Z(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09118_ (.A1(_02353_),
    .A2(_03518_),
    .ZN(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09119_ (.I(_03505_),
    .ZN(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _09120_ (.A1(_03506_),
    .A2(_03492_),
    .B(_03521_),
    .C(_03507_),
    .ZN(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09121_ (.A1(_03520_),
    .A2(_03522_),
    .ZN(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09122_ (.A1(_02367_),
    .A2(_03519_),
    .A3(_03523_),
    .Z(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09123_ (.A1(_03471_),
    .A2(_03524_),
    .B(_03510_),
    .ZN(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09124_ (.A1(_03516_),
    .A2(_03502_),
    .B1(_03525_),
    .B2(_01666_),
    .ZN(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09125_ (.A1(\as2650.instruction_args_latch[7] ),
    .A2(_03397_),
    .ZN(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09126_ (.A1(_01669_),
    .A2(_03398_),
    .B(_03527_),
    .ZN(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09127_ (.A1(_03468_),
    .A2(_03526_),
    .B1(_03528_),
    .B2(_03394_),
    .ZN(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09128_ (.A1(_03516_),
    .A2(_03467_),
    .B(_03517_),
    .C(_03529_),
    .ZN(_00383_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09129_ (.I(\as2650.indirect_target[8] ),
    .ZN(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09130_ (.A1(_02383_),
    .A2(_03518_),
    .ZN(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09131_ (.A1(_02382_),
    .A2(_03518_),
    .Z(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09132_ (.A1(_03531_),
    .A2(_03532_),
    .ZN(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09133_ (.I(_03504_),
    .Z(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09134_ (.A1(_02367_),
    .A2(_03534_),
    .ZN(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09135_ (.A1(_02367_),
    .A2(_03534_),
    .ZN(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _09136_ (.A1(_03522_),
    .A2(_03535_),
    .B(_03536_),
    .C(_03520_),
    .ZN(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09137_ (.A1(_03533_),
    .A2(_03537_),
    .ZN(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09138_ (.A1(_03381_),
    .A2(_03538_),
    .B(_03510_),
    .ZN(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09139_ (.A1(_03530_),
    .A2(_03502_),
    .B1(_03539_),
    .B2(_01666_),
    .ZN(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09140_ (.I(_03375_),
    .Z(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09141_ (.A1(_03385_),
    .A2(_03423_),
    .B1(_03540_),
    .B2(_03541_),
    .ZN(_03542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09142_ (.A1(_03530_),
    .A2(_01440_),
    .B(_03517_),
    .C(_03542_),
    .ZN(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09143_ (.I(_01354_),
    .Z(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09144_ (.I(_03543_),
    .Z(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09145_ (.I(_01348_),
    .Z(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09146_ (.A1(_03373_),
    .A2(_03374_),
    .A3(_02875_),
    .ZN(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09147_ (.I(_03546_),
    .Z(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09148_ (.I(_03388_),
    .Z(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09149_ (.A1(_02398_),
    .A2(_03504_),
    .ZN(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09150_ (.A1(_02383_),
    .A2(_03534_),
    .Z(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09151_ (.A1(_03532_),
    .A2(_03537_),
    .B(_03550_),
    .ZN(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09152_ (.A1(_03549_),
    .A2(_03551_),
    .Z(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09153_ (.I(net296),
    .ZN(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09154_ (.A1(_03553_),
    .A2(_03381_),
    .ZN(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09155_ (.I(_03554_),
    .Z(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09156_ (.A1(\as2650.indirect_target[9] ),
    .A2(_03548_),
    .B1(_03552_),
    .B2(_03555_),
    .ZN(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09157_ (.A1(_03541_),
    .A2(_03556_),
    .ZN(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09158_ (.A1(\as2650.indirect_target[9] ),
    .A2(_03545_),
    .B1(_03547_),
    .B2(_03408_),
    .C(_03557_),
    .ZN(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09159_ (.A1(_03544_),
    .A2(_03558_),
    .ZN(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09160_ (.I(_03546_),
    .Z(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09161_ (.A1(_02412_),
    .A2(_03519_),
    .ZN(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09162_ (.I(_03534_),
    .Z(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09163_ (.A1(_03533_),
    .A2(_03549_),
    .ZN(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09164_ (.A1(_02398_),
    .A2(_03561_),
    .B1(_03537_),
    .B2(_03562_),
    .C(_03550_),
    .ZN(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09165_ (.A1(_03560_),
    .A2(_03563_),
    .ZN(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09166_ (.A1(\as2650.indirect_target[10] ),
    .A2(_03548_),
    .ZN(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09167_ (.A1(_03553_),
    .A2(_03471_),
    .A3(_03564_),
    .B(_03565_),
    .ZN(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09168_ (.I(_03541_),
    .ZN(_03567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _09169_ (.A1(\as2650.indirect_target[10] ),
    .A2(_03545_),
    .B1(_03559_),
    .B2(_03428_),
    .C1(_03566_),
    .C2(_03567_),
    .ZN(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09170_ (.A1(_03544_),
    .A2(_03568_),
    .ZN(_00386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09171_ (.A1(\as2650.instruction_args_latch[11] ),
    .A2(_03486_),
    .ZN(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09172_ (.A1(_03452_),
    .A2(_03486_),
    .B(_03569_),
    .ZN(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09173_ (.I(_03570_),
    .Z(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09174_ (.A1(_02421_),
    .A2(_03519_),
    .ZN(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09175_ (.I(_02412_),
    .Z(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09176_ (.A1(_03573_),
    .A2(_03561_),
    .ZN(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09177_ (.A1(_03573_),
    .A2(_03561_),
    .ZN(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09178_ (.A1(_03574_),
    .A2(_03563_),
    .B(_03575_),
    .ZN(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09179_ (.A1(_03572_),
    .A2(_03576_),
    .ZN(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09180_ (.A1(\as2650.indirect_target[11] ),
    .A2(_03548_),
    .B1(_03554_),
    .B2(_03577_),
    .ZN(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09181_ (.A1(_03541_),
    .A2(_03578_),
    .ZN(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09182_ (.A1(\as2650.indirect_target[11] ),
    .A2(_03545_),
    .B1(_03547_),
    .B2(_03571_),
    .C(_03579_),
    .ZN(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09183_ (.A1(_03544_),
    .A2(_03580_),
    .ZN(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09184_ (.I(_03519_),
    .Z(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09185_ (.A1(_02413_),
    .A2(_02421_),
    .B(_03561_),
    .ZN(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09186_ (.A1(_03560_),
    .A2(_03563_),
    .A3(_03572_),
    .B(_03582_),
    .ZN(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09187_ (.A1(_02441_),
    .A2(_03581_),
    .A3(_03583_),
    .Z(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09188_ (.A1(\as2650.indirect_target[12] ),
    .A2(_03548_),
    .B1(_03554_),
    .B2(_03584_),
    .ZN(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09189_ (.A1(_03375_),
    .A2(_03585_),
    .ZN(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09190_ (.A1(\as2650.indirect_target[12] ),
    .A2(_03545_),
    .B1(_03547_),
    .B2(_03490_),
    .C(_03586_),
    .ZN(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09191_ (.A1(_03544_),
    .A2(_03587_),
    .ZN(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09192_ (.I(_01448_),
    .Z(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09193_ (.A1(\as2650.indirect_target[13] ),
    .A2(_03389_),
    .B1(_03555_),
    .B2(_02448_),
    .ZN(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09194_ (.I(_00722_),
    .Z(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09195_ (.I(_03488_),
    .Z(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09196_ (.A1(_02145_),
    .A2(_03591_),
    .Z(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09197_ (.A1(_02448_),
    .A2(_03590_),
    .B(_03559_),
    .C(_03592_),
    .ZN(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09198_ (.A1(_03547_),
    .A2(_03589_),
    .B(_03593_),
    .ZN(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09199_ (.A1(_03588_),
    .A2(_03594_),
    .Z(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09200_ (.I(_03595_),
    .Z(_00389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09201_ (.I(_03543_),
    .Z(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09202_ (.I(_03546_),
    .Z(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09203_ (.I0(_02457_),
    .I1(_03581_),
    .S(_03590_),
    .Z(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09204_ (.A1(\as2650.indirect_target[14] ),
    .A2(_03502_),
    .B1(_03555_),
    .B2(_02457_),
    .ZN(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09205_ (.A1(_03559_),
    .A2(_03599_),
    .ZN(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09206_ (.A1(_03597_),
    .A2(_03598_),
    .B(_03600_),
    .ZN(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09207_ (.A1(_03596_),
    .A2(_03601_),
    .ZN(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09208_ (.A1(_03597_),
    .A2(_03555_),
    .B(_02466_),
    .ZN(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09209_ (.A1(\as2650.indirect_target[15] ),
    .A2(_03389_),
    .A3(_03423_),
    .ZN(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09210_ (.I(_01684_),
    .Z(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09211_ (.A1(_03602_),
    .A2(_03603_),
    .B(_03604_),
    .ZN(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09212_ (.I(_00908_),
    .ZN(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09213_ (.I(_02258_),
    .Z(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09214_ (.A1(_03606_),
    .A2(_03559_),
    .ZN(_03607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09215_ (.A1(_03605_),
    .A2(_03597_),
    .B1(_03607_),
    .B2(\as2650.indexed_cyc[0] ),
    .ZN(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09216_ (.A1(_01448_),
    .A2(_02961_),
    .ZN(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09217_ (.I(_03609_),
    .Z(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09218_ (.A1(_03608_),
    .A2(_03610_),
    .ZN(_00392_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09219_ (.I(_00734_),
    .ZN(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09220_ (.A1(_03611_),
    .A2(_03597_),
    .B1(_03607_),
    .B2(\as2650.indexed_cyc[1] ),
    .ZN(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09221_ (.A1(_03610_),
    .A2(_03612_),
    .ZN(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09222_ (.I(_02149_),
    .Z(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09223_ (.I(_01387_),
    .Z(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09224_ (.A1(_03373_),
    .A2(_01664_),
    .ZN(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09225_ (.A1(_00925_),
    .A2(_03613_),
    .B1(_03614_),
    .B2(_03615_),
    .ZN(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09226_ (.A1(_03466_),
    .A2(_03616_),
    .ZN(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09227_ (.A1(_00658_),
    .A2(_01514_),
    .B1(_03393_),
    .B2(_03617_),
    .ZN(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09228_ (.A1(_03610_),
    .A2(_03618_),
    .ZN(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09229_ (.I(_01683_),
    .Z(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09230_ (.I(_03619_),
    .Z(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09231_ (.A1(_02258_),
    .A2(_01654_),
    .ZN(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09232_ (.I(_03621_),
    .Z(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09233_ (.A1(_03622_),
    .A2(_02866_),
    .ZN(_03623_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09234_ (.A1(net196),
    .A2(_03623_),
    .ZN(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09235_ (.A1(_01268_),
    .A2(_01655_),
    .Z(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09236_ (.A1(_03620_),
    .A2(_03624_),
    .A3(_03625_),
    .ZN(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09237_ (.A1(_03613_),
    .A2(_02873_),
    .B(_01187_),
    .ZN(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09238_ (.A1(_02864_),
    .A2(_02147_),
    .B(_03614_),
    .ZN(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09239_ (.A1(_03626_),
    .A2(_03627_),
    .B(_03369_),
    .ZN(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09240_ (.I(_01520_),
    .Z(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09241_ (.I(_03629_),
    .Z(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09242_ (.I(_03630_),
    .Z(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09243_ (.I(_03631_),
    .Z(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09244_ (.I(_02846_),
    .Z(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09245_ (.A1(_03411_),
    .A2(_03633_),
    .A3(_01507_),
    .A4(_02841_),
    .ZN(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09246_ (.A1(_01503_),
    .A2(_01442_),
    .A3(_02833_),
    .A4(_02156_),
    .ZN(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09247_ (.A1(_02834_),
    .A2(_03635_),
    .ZN(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09248_ (.A1(_01504_),
    .A2(_02201_),
    .A3(_01376_),
    .ZN(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09249_ (.A1(_02843_),
    .A2(_03634_),
    .A3(_03636_),
    .A4(_03637_),
    .Z(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09250_ (.A1(_01660_),
    .A2(_03638_),
    .ZN(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09251_ (.I(_03639_),
    .Z(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09252_ (.I(_03640_),
    .Z(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09253_ (.A1(_03632_),
    .A2(_03641_),
    .B(_02229_),
    .ZN(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09254_ (.I(_03629_),
    .Z(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09255_ (.I(_03643_),
    .Z(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09256_ (.I(_03644_),
    .Z(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09257_ (.A1(_03645_),
    .A2(_03634_),
    .A3(_03641_),
    .Z(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09258_ (.A1(_03517_),
    .A2(_03628_),
    .A3(_03642_),
    .A4(_03646_),
    .ZN(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09259_ (.I(_03647_),
    .Z(_00396_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09260_ (.I(\as2650.warmup[1] ),
    .ZN(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09261_ (.A1(\as2650.warmup[0] ),
    .A2(_03648_),
    .B(_01252_),
    .ZN(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09262_ (.A1(\as2650.warmup[0] ),
    .A2(\as2650.warmup[1] ),
    .ZN(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09263_ (.A1(_01252_),
    .A2(_03649_),
    .ZN(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09264_ (.I(_03392_),
    .Z(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09265_ (.I(_03650_),
    .Z(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09266_ (.I(_03392_),
    .Z(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09267_ (.A1(_03606_),
    .A2(_03652_),
    .ZN(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09268_ (.I(_03653_),
    .Z(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09269_ (.A1(_02892_),
    .A2(_03651_),
    .B1(_03654_),
    .B2(\as2650.instruction_args_latch[0] ),
    .ZN(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09270_ (.A1(_03610_),
    .A2(_03655_),
    .ZN(_00399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09271_ (.I(_03609_),
    .Z(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09272_ (.I(_03656_),
    .Z(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09273_ (.I(_03406_),
    .Z(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09274_ (.A1(_03658_),
    .A2(_03651_),
    .B1(_03654_),
    .B2(\as2650.instruction_args_latch[1] ),
    .ZN(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09275_ (.A1(_03657_),
    .A2(_03659_),
    .ZN(_00400_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09276_ (.I(_03433_),
    .Z(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09277_ (.A1(_03660_),
    .A2(_03651_),
    .B1(_03654_),
    .B2(\as2650.instruction_args_latch[2] ),
    .ZN(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09278_ (.A1(_03657_),
    .A2(_03661_),
    .ZN(_00401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09279_ (.A1(_03094_),
    .A2(_03651_),
    .B1(_03654_),
    .B2(\as2650.instruction_args_latch[3] ),
    .ZN(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09280_ (.A1(_03657_),
    .A2(_03662_),
    .ZN(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09281_ (.I(_03470_),
    .Z(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09282_ (.I(_03652_),
    .Z(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09283_ (.I(_03653_),
    .Z(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09284_ (.A1(_03663_),
    .A2(_03664_),
    .B1(_03665_),
    .B2(\as2650.instruction_args_latch[4] ),
    .ZN(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09285_ (.A1(_03657_),
    .A2(_03666_),
    .ZN(_00403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09286_ (.A1(_00695_),
    .A2(net123),
    .B(_00696_),
    .ZN(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09287_ (.I(_03667_),
    .Z(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09288_ (.I(_03668_),
    .Z(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09289_ (.A1(_03669_),
    .A2(_03664_),
    .B1(_03665_),
    .B2(\as2650.instruction_args_latch[5] ),
    .ZN(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09290_ (.A1(_03656_),
    .A2(_03670_),
    .ZN(_00404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09291_ (.I(_03243_),
    .Z(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09292_ (.I(_03671_),
    .Z(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09293_ (.A1(_03672_),
    .A2(_03664_),
    .B1(_03665_),
    .B2(\as2650.instruction_args_latch[6] ),
    .ZN(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09294_ (.A1(_03656_),
    .A2(_03673_),
    .ZN(_00405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09295_ (.A1(_00701_),
    .A2(net123),
    .B(_00702_),
    .ZN(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09296_ (.I(_03674_),
    .Z(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09297_ (.A1(_03675_),
    .A2(_03664_),
    .B1(_03665_),
    .B2(\as2650.instruction_args_latch[7] ),
    .ZN(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09298_ (.A1(_03656_),
    .A2(_03676_),
    .ZN(_00406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09299_ (.I(_02960_),
    .Z(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09300_ (.I(_03677_),
    .Z(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09301_ (.I(_02863_),
    .Z(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _09302_ (.A1(_03679_),
    .A2(_03625_),
    .Z(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09303_ (.A1(_03606_),
    .A2(_03678_),
    .A3(_03680_),
    .ZN(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09304_ (.I(_03681_),
    .Z(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09305_ (.A1(\as2650.instruction_args_latch[8] ),
    .A2(_03682_),
    .ZN(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09306_ (.I(_03680_),
    .Z(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09307_ (.A1(_02892_),
    .A2(_03684_),
    .ZN(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09308_ (.A1(_03683_),
    .A2(_03685_),
    .B(_03604_),
    .ZN(_00407_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09309_ (.A1(_03658_),
    .A2(_03684_),
    .B1(_03682_),
    .B2(\as2650.instruction_args_latch[9] ),
    .ZN(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09310_ (.A1(_03596_),
    .A2(_03686_),
    .ZN(_00408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09311_ (.A1(_03660_),
    .A2(_03684_),
    .B1(_03682_),
    .B2(\as2650.instruction_args_latch[10] ),
    .ZN(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09312_ (.A1(_03596_),
    .A2(_03687_),
    .ZN(_00409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09313_ (.A1(_03094_),
    .A2(_03684_),
    .B1(_03682_),
    .B2(\as2650.instruction_args_latch[11] ),
    .ZN(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09314_ (.A1(_03596_),
    .A2(_03688_),
    .ZN(_00410_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09315_ (.I(_03543_),
    .Z(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09316_ (.I(_03680_),
    .Z(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09317_ (.I(_03681_),
    .Z(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09318_ (.A1(_03663_),
    .A2(_03690_),
    .B1(_03691_),
    .B2(\as2650.instruction_args_latch[12] ),
    .ZN(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09319_ (.A1(_03689_),
    .A2(_03692_),
    .ZN(_00411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09320_ (.A1(_03669_),
    .A2(_03690_),
    .B1(_03691_),
    .B2(_00723_),
    .ZN(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09321_ (.A1(_03689_),
    .A2(_03693_),
    .ZN(_00412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09322_ (.A1(_03672_),
    .A2(_03690_),
    .B1(_03691_),
    .B2(\as2650.instruction_args_latch[14] ),
    .ZN(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09323_ (.A1(_03689_),
    .A2(_03694_),
    .ZN(_00413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09324_ (.A1(_03675_),
    .A2(_03690_),
    .B1(_03691_),
    .B2(\as2650.instruction_args_latch[15] ),
    .ZN(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09325_ (.A1(_03689_),
    .A2(_03695_),
    .ZN(_00414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09326_ (.I(_02152_),
    .Z(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09327_ (.I(_03630_),
    .Z(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09328_ (.A1(_01664_),
    .A2(_02146_),
    .B(_03614_),
    .ZN(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09329_ (.I(_02830_),
    .Z(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09330_ (.I(_03699_),
    .Z(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09331_ (.I(_02866_),
    .ZN(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09332_ (.A1(_01660_),
    .A2(_03701_),
    .A3(_03638_),
    .ZN(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09333_ (.A1(_03700_),
    .A2(_03702_),
    .B(_03606_),
    .ZN(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09334_ (.A1(_03626_),
    .A2(_03698_),
    .A3(_03703_),
    .Z(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09335_ (.A1(_03696_),
    .A2(_03697_),
    .A3(_03650_),
    .B1(_03704_),
    .B2(_03466_),
    .ZN(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09336_ (.I(_02856_),
    .Z(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09337_ (.A1(_01356_),
    .A2(_01361_),
    .B(_03706_),
    .C(_03625_),
    .ZN(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09338_ (.A1(_01361_),
    .A2(_03705_),
    .B(_03707_),
    .ZN(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09339_ (.A1(net40),
    .A2(net39),
    .A3(net41),
    .ZN(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09340_ (.A1(net36),
    .A2(net35),
    .A3(net38),
    .A4(net37),
    .ZN(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09341_ (.A1(_01360_),
    .A2(_00931_),
    .ZN(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09342_ (.A1(_02258_),
    .A2(_01346_),
    .B1(_03711_),
    .B2(_02855_),
    .ZN(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09343_ (.A1(_03709_),
    .A2(_03710_),
    .B(_01896_),
    .C(_03712_),
    .ZN(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09344_ (.I(_03713_),
    .ZN(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09345_ (.A1(_03696_),
    .A2(_03706_),
    .ZN(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09346_ (.A1(_01347_),
    .A2(_02154_),
    .ZN(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09347_ (.I(_03716_),
    .Z(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09348_ (.A1(_03440_),
    .A2(_03717_),
    .ZN(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09349_ (.A1(_03708_),
    .A2(_03714_),
    .A3(_03715_),
    .A4(_03718_),
    .Z(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09350_ (.I(_03719_),
    .Z(_00415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09351_ (.I(_01385_),
    .Z(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09352_ (.I(_02875_),
    .Z(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09353_ (.I(_01679_),
    .Z(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09354_ (.A1(_03722_),
    .A2(_01661_),
    .B(_00645_),
    .ZN(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09355_ (.A1(_03623_),
    .A2(_03723_),
    .B(_03627_),
    .ZN(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _09356_ (.A1(_03590_),
    .A2(_03721_),
    .A3(_03393_),
    .B1(_03724_),
    .B2(_03613_),
    .ZN(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _09357_ (.A1(_03720_),
    .A2(_03369_),
    .B1(_03706_),
    .B2(_00931_),
    .C1(_03725_),
    .C2(_01224_),
    .ZN(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09358_ (.A1(_01433_),
    .A2(_02857_),
    .ZN(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09359_ (.A1(_03696_),
    .A2(_03720_),
    .A3(_02855_),
    .A4(_01244_),
    .ZN(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09360_ (.I(_03728_),
    .Z(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09361_ (.A1(_03727_),
    .A2(_03729_),
    .ZN(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09362_ (.A1(_01179_),
    .A2(_01440_),
    .B(_03714_),
    .C(_03730_),
    .ZN(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09363_ (.A1(_03726_),
    .A2(_03731_),
    .ZN(_00416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09364_ (.A1(_01360_),
    .A2(_03466_),
    .B(_03720_),
    .ZN(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09365_ (.A1(_01382_),
    .A2(_03701_),
    .B(_01244_),
    .ZN(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09366_ (.A1(_03720_),
    .A2(_01348_),
    .A3(_03733_),
    .ZN(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09367_ (.A1(_02855_),
    .A2(_03734_),
    .ZN(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09368_ (.A1(_00934_),
    .A2(_03732_),
    .B1(_03735_),
    .B2(_03696_),
    .C(_03714_),
    .ZN(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09369_ (.A1(_03588_),
    .A2(_03736_),
    .Z(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09370_ (.I(_03737_),
    .Z(_00417_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _09371_ (.A1(_01505_),
    .A2(_02833_),
    .ZN(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09372_ (.I(_00788_),
    .Z(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _09373_ (.A1(_03739_),
    .A2(_03255_),
    .A3(_02842_),
    .ZN(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09374_ (.A1(_01411_),
    .A2(_03740_),
    .ZN(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09375_ (.A1(_01679_),
    .A2(_01663_),
    .A3(_03741_),
    .ZN(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09376_ (.A1(_01462_),
    .A2(_01509_),
    .A3(_03738_),
    .A4(_03742_),
    .Z(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09377_ (.I(_03743_),
    .Z(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09378_ (.A1(_02152_),
    .A2(_02153_),
    .A3(_01655_),
    .ZN(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09379_ (.I(_03745_),
    .Z(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09380_ (.I(_03746_),
    .Z(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09381_ (.A1(_01360_),
    .A2(_03744_),
    .B(_03747_),
    .C(_02857_),
    .ZN(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09382_ (.A1(_03625_),
    .A2(_03713_),
    .ZN(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09383_ (.A1(_03748_),
    .A2(_03749_),
    .B(_03604_),
    .ZN(_00418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09384_ (.A1(net30),
    .A2(_03180_),
    .B(_00740_),
    .ZN(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09385_ (.I(_03750_),
    .Z(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09386_ (.I(_03751_),
    .Z(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09387_ (.I(_03644_),
    .Z(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09388_ (.I(_03753_),
    .Z(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09389_ (.A1(\as2650.insin[0] ),
    .A2(_03632_),
    .ZN(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09390_ (.I(_03619_),
    .Z(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09391_ (.A1(_03752_),
    .A2(_03754_),
    .B(_03755_),
    .C(_03756_),
    .ZN(_00419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09392_ (.I(_02977_),
    .Z(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09393_ (.A1(\as2650.insin[1] ),
    .A2(_03632_),
    .ZN(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09394_ (.I(_03440_),
    .Z(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09395_ (.A1(_03757_),
    .A2(_03754_),
    .B(_03758_),
    .C(_03759_),
    .ZN(_00420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09396_ (.I(_03042_),
    .Z(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09397_ (.A1(\as2650.insin[2] ),
    .A2(_03632_),
    .ZN(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09398_ (.A1(_03760_),
    .A2(_03754_),
    .B(_03761_),
    .C(_03759_),
    .ZN(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09399_ (.I(_03453_),
    .Z(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09400_ (.I(_03697_),
    .Z(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09401_ (.A1(\as2650.insin[3] ),
    .A2(_03763_),
    .ZN(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09402_ (.A1(_03762_),
    .A2(_03754_),
    .B(_03764_),
    .C(_03759_),
    .ZN(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09403_ (.I(_03182_),
    .Z(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09404_ (.I(_03753_),
    .Z(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09405_ (.A1(\as2650.insin[4] ),
    .A2(_03763_),
    .ZN(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09406_ (.A1(_03765_),
    .A2(_03766_),
    .B(_03767_),
    .C(_03759_),
    .ZN(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09407_ (.I(_03196_),
    .Z(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09408_ (.A1(\as2650.insin[5] ),
    .A2(_03763_),
    .ZN(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09409_ (.I(_03440_),
    .Z(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09410_ (.A1(_03768_),
    .A2(_03766_),
    .B(_03769_),
    .C(_03770_),
    .ZN(_00424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09411_ (.I(_03241_),
    .Z(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09412_ (.A1(\as2650.insin[6] ),
    .A2(_03763_),
    .ZN(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09413_ (.A1(_03771_),
    .A2(_03766_),
    .B(_03772_),
    .C(_03770_),
    .ZN(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09414_ (.I(_03291_),
    .Z(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09415_ (.A1(\as2650.insin[7] ),
    .A2(_03753_),
    .ZN(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09416_ (.A1(_03773_),
    .A2(_03766_),
    .B(_03774_),
    .C(_03770_),
    .ZN(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09417_ (.I(_03543_),
    .Z(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09418_ (.I(_03746_),
    .Z(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _09419_ (.A1(_03383_),
    .A2(_03384_),
    .Z(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09420_ (.I(_03428_),
    .ZN(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09421_ (.I(_02204_),
    .Z(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09422_ (.A1(net195),
    .A2(_03779_),
    .ZN(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _09423_ (.A1(_03528_),
    .A2(_03780_),
    .ZN(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09424_ (.I(_03779_),
    .Z(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09425_ (.A1(net194),
    .A2(_03782_),
    .B(_03514_),
    .ZN(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09426_ (.A1(net192),
    .A2(_02205_),
    .ZN(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _09427_ (.A1(_03499_),
    .A2(_03784_),
    .ZN(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09428_ (.A1(net191),
    .A2(_03779_),
    .B(_03482_),
    .ZN(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09429_ (.A1(net190),
    .A2(_02204_),
    .ZN(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _09430_ (.A1(_03462_),
    .A2(_03787_),
    .ZN(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09431_ (.A1(net189),
    .A2(_02204_),
    .B(_03437_),
    .ZN(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09432_ (.A1(net188),
    .A2(_02203_),
    .ZN(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09433_ (.A1(_03420_),
    .A2(_03421_),
    .A3(_03790_),
    .ZN(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09434_ (.A1(net187),
    .A2(_02203_),
    .ZN(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09435_ (.A1(_01008_),
    .A2(_03396_),
    .B(_03399_),
    .C(_03792_),
    .ZN(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09436_ (.A1(_03420_),
    .A2(_03421_),
    .B(_03790_),
    .ZN(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09437_ (.A1(_03791_),
    .A2(_03793_),
    .B(_03794_),
    .ZN(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09438_ (.A1(net189),
    .A2(_02205_),
    .A3(_03437_),
    .ZN(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09439_ (.A1(_03789_),
    .A2(_03795_),
    .B(_03796_),
    .ZN(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09440_ (.A1(net190),
    .A2(_02205_),
    .A3(_03462_),
    .Z(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09441_ (.A1(_03788_),
    .A2(_03797_),
    .B(_03798_),
    .ZN(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09442_ (.A1(net191),
    .A2(_03779_),
    .A3(_03482_),
    .ZN(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09443_ (.A1(_03786_),
    .A2(_03799_),
    .B(_03800_),
    .ZN(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09444_ (.A1(net192),
    .A2(_03782_),
    .A3(_03499_),
    .Z(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09445_ (.A1(_03785_),
    .A2(_03801_),
    .B(_03802_),
    .ZN(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09446_ (.A1(net194),
    .A2(_03782_),
    .A3(_03514_),
    .ZN(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09447_ (.A1(_03783_),
    .A2(_03803_),
    .B(_03804_),
    .ZN(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09448_ (.I(_03782_),
    .Z(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09449_ (.A1(net195),
    .A2(_03806_),
    .A3(_03528_),
    .Z(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09450_ (.A1(_03781_),
    .A2(_03805_),
    .B(_03807_),
    .ZN(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09451_ (.A1(_03777_),
    .A2(_03409_),
    .A3(_03778_),
    .A4(_03808_),
    .ZN(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09452_ (.A1(_03570_),
    .A2(_03490_),
    .A3(_03809_),
    .Z(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09453_ (.A1(_02873_),
    .A2(_02210_),
    .Z(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09454_ (.I(_03811_),
    .Z(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09455_ (.A1(_03391_),
    .A2(_03812_),
    .Z(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09456_ (.I(_03813_),
    .Z(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09457_ (.A1(_03591_),
    .A2(_03810_),
    .B(_03814_),
    .ZN(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09458_ (.A1(_03591_),
    .A2(_03810_),
    .Z(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09459_ (.I(_03746_),
    .Z(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09460_ (.A1(_03391_),
    .A2(_03812_),
    .ZN(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09461_ (.A1(_02198_),
    .A2(_03738_),
    .Z(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09462_ (.I(_03819_),
    .Z(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09463_ (.A1(_03629_),
    .A2(_03820_),
    .ZN(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09464_ (.A1(\as2650.debug_psu[3] ),
    .A2(_02533_),
    .Z(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09465_ (.I(_03822_),
    .Z(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09466_ (.I(_03823_),
    .Z(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09467_ (.I(_03824_),
    .Z(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09468_ (.I(_03825_),
    .Z(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _09469_ (.A1(\as2650.debug_psu[0] ),
    .A2(_01858_),
    .ZN(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09470_ (.A1(_02246_),
    .A2(_03827_),
    .Z(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09471_ (.I(_03828_),
    .Z(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09472_ (.I(_03829_),
    .Z(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09473_ (.I(_03830_),
    .Z(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09474_ (.I(_02253_),
    .Z(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09475_ (.I(_03827_),
    .Z(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09476_ (.I(_03833_),
    .Z(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09477_ (.I(_03834_),
    .Z(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09478_ (.I(_03835_),
    .Z(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09479_ (.I(_03836_),
    .Z(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09480_ (.A1(\as2650.stack[10][13] ),
    .A2(_03832_),
    .B1(_03837_),
    .B2(\as2650.stack[11][13] ),
    .ZN(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09481_ (.I(_02480_),
    .Z(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09482_ (.I(_02597_),
    .Z(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09483_ (.A1(\as2650.stack[9][13] ),
    .A2(_03839_),
    .B1(_03840_),
    .B2(\as2650.stack[8][13] ),
    .ZN(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09484_ (.A1(_03831_),
    .A2(_03838_),
    .A3(_03841_),
    .ZN(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09485_ (.A1(\as2650.debug_psu[2] ),
    .A2(_03827_),
    .Z(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09486_ (.I(_03843_),
    .Z(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09487_ (.I(_03844_),
    .Z(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09488_ (.I(_03845_),
    .Z(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09489_ (.I(_03846_),
    .Z(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09490_ (.I(_02480_),
    .Z(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09491_ (.I(_02597_),
    .Z(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09492_ (.A1(\as2650.stack[13][13] ),
    .A2(_03848_),
    .B1(_03849_),
    .B2(\as2650.stack[12][13] ),
    .ZN(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09493_ (.I(_02253_),
    .Z(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09494_ (.I(_03836_),
    .Z(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09495_ (.A1(\as2650.stack[14][13] ),
    .A2(_03851_),
    .B1(_03852_),
    .B2(\as2650.stack[15][13] ),
    .ZN(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09496_ (.A1(_03847_),
    .A2(_03850_),
    .A3(_03853_),
    .ZN(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09497_ (.A1(_03842_),
    .A2(_03854_),
    .Z(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09498_ (.I(_02253_),
    .Z(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09499_ (.I(_03836_),
    .Z(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09500_ (.A1(\as2650.stack[5][13] ),
    .A2(_02480_),
    .B1(_02597_),
    .B2(\as2650.stack[4][13] ),
    .ZN(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09501_ (.I(_03858_),
    .ZN(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09502_ (.A1(\as2650.stack[6][13] ),
    .A2(_03856_),
    .B1(_03857_),
    .B2(\as2650.stack[7][13] ),
    .C(_03859_),
    .ZN(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09503_ (.A1(_03847_),
    .A2(_03860_),
    .B(_03825_),
    .ZN(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09504_ (.I(_03831_),
    .Z(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09505_ (.A1(\as2650.stack[2][13] ),
    .A2(_02254_),
    .B1(_03857_),
    .B2(\as2650.stack[3][13] ),
    .ZN(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09506_ (.A1(\as2650.stack[1][13] ),
    .A2(_02481_),
    .B1(_02598_),
    .B2(\as2650.stack[0][13] ),
    .ZN(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09507_ (.A1(_03862_),
    .A2(_03863_),
    .A3(_03864_),
    .ZN(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _09508_ (.A1(_03826_),
    .A2(_03855_),
    .B1(_03861_),
    .B2(_03865_),
    .ZN(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09509_ (.A1(_03615_),
    .A2(_03811_),
    .Z(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09510_ (.I(_03867_),
    .Z(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09511_ (.A1(_03679_),
    .A2(_03868_),
    .ZN(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09512_ (.A1(_03377_),
    .A2(_03869_),
    .B(_03821_),
    .C(_02448_),
    .ZN(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09513_ (.A1(_03821_),
    .A2(_03866_),
    .B(_03870_),
    .ZN(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09514_ (.A1(_03818_),
    .A2(_03871_),
    .ZN(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09515_ (.A1(_03815_),
    .A2(_03816_),
    .B(_03817_),
    .C(_03872_),
    .ZN(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09516_ (.A1(_00723_),
    .A2(_03776_),
    .B(_03873_),
    .ZN(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09517_ (.A1(_03775_),
    .A2(_03874_),
    .ZN(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09518_ (.I(_03717_),
    .Z(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09519_ (.I(_03813_),
    .Z(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09520_ (.I(_03876_),
    .Z(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09521_ (.A1(_03581_),
    .A2(_03816_),
    .Z(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09522_ (.I(_03876_),
    .Z(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09523_ (.A1(_03377_),
    .A2(_03868_),
    .ZN(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09524_ (.A1(_03722_),
    .A2(_03880_),
    .ZN(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09525_ (.A1(\as2650.stack[2][14] ),
    .A2(_03832_),
    .B1(_03852_),
    .B2(\as2650.stack[3][14] ),
    .ZN(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09526_ (.A1(\as2650.stack[1][14] ),
    .A2(_03848_),
    .B1(_03849_),
    .B2(\as2650.stack[0][14] ),
    .ZN(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09527_ (.A1(_03831_),
    .A2(_03882_),
    .A3(_03883_),
    .ZN(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09528_ (.A1(\as2650.stack[5][14] ),
    .A2(_03839_),
    .B1(_03840_),
    .B2(\as2650.stack[4][14] ),
    .ZN(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09529_ (.A1(\as2650.stack[6][14] ),
    .A2(_03851_),
    .B1(_03852_),
    .B2(\as2650.stack[7][14] ),
    .ZN(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09530_ (.A1(_03846_),
    .A2(_03885_),
    .A3(_03886_),
    .ZN(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09531_ (.A1(_03884_),
    .A2(_03887_),
    .ZN(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09532_ (.A1(\as2650.stack[10][14] ),
    .A2(_03851_),
    .B1(_03852_),
    .B2(\as2650.stack[11][14] ),
    .ZN(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09533_ (.A1(\as2650.stack[9][14] ),
    .A2(_03839_),
    .B1(_03840_),
    .B2(\as2650.stack[8][14] ),
    .ZN(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09534_ (.A1(_03831_),
    .A2(_03889_),
    .A3(_03890_),
    .ZN(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09535_ (.A1(\as2650.stack[13][14] ),
    .A2(_03839_),
    .B1(_03840_),
    .B2(\as2650.stack[12][14] ),
    .ZN(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09536_ (.A1(\as2650.stack[14][14] ),
    .A2(_03851_),
    .B1(_03836_),
    .B2(\as2650.stack[15][14] ),
    .ZN(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09537_ (.A1(_03846_),
    .A2(_03892_),
    .A3(_03893_),
    .ZN(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09538_ (.A1(_03825_),
    .A2(_03891_),
    .A3(_03894_),
    .ZN(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09539_ (.A1(_03826_),
    .A2(_03888_),
    .B(_03895_),
    .ZN(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09540_ (.I0(_03896_),
    .I1(\as2650.page_reg[1] ),
    .S(_03821_),
    .Z(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09541_ (.A1(_02457_),
    .A2(_03881_),
    .B1(_03897_),
    .B2(_03869_),
    .ZN(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09542_ (.I(_03745_),
    .Z(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09543_ (.A1(_03879_),
    .A2(_03898_),
    .B(_03899_),
    .ZN(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09544_ (.A1(_03877_),
    .A2(_03878_),
    .B(_03900_),
    .ZN(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09545_ (.A1(_00731_),
    .A2(_03875_),
    .B(_03901_),
    .C(_03770_),
    .ZN(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09546_ (.A1(_03591_),
    .A2(_03581_),
    .A3(_03810_),
    .ZN(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09547_ (.I0(_01673_),
    .I1(\as2650.page_reg[2] ),
    .S(_01228_),
    .Z(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09548_ (.A1(_03902_),
    .A2(_03903_),
    .ZN(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09549_ (.A1(\as2650.stack[2][15] ),
    .A2(_03856_),
    .B1(_03857_),
    .B2(\as2650.stack[3][15] ),
    .ZN(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09550_ (.A1(\as2650.stack[1][15] ),
    .A2(_02481_),
    .B1(_02598_),
    .B2(\as2650.stack[0][15] ),
    .ZN(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09551_ (.A1(_03862_),
    .A2(_03905_),
    .A3(_03906_),
    .ZN(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09552_ (.A1(\as2650.stack[5][15] ),
    .A2(_02481_),
    .B1(_02598_),
    .B2(\as2650.stack[4][15] ),
    .ZN(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09553_ (.A1(\as2650.stack[6][15] ),
    .A2(_03856_),
    .B1(_03837_),
    .B2(\as2650.stack[7][15] ),
    .ZN(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09554_ (.A1(_03847_),
    .A2(_03908_),
    .A3(_03909_),
    .ZN(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09555_ (.A1(_03907_),
    .A2(_03910_),
    .ZN(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09556_ (.A1(\as2650.stack[10][15] ),
    .A2(_03832_),
    .B1(_03837_),
    .B2(\as2650.stack[11][15] ),
    .ZN(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09557_ (.A1(\as2650.stack[9][15] ),
    .A2(_03848_),
    .B1(_03849_),
    .B2(\as2650.stack[8][15] ),
    .ZN(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09558_ (.A1(_03862_),
    .A2(_03912_),
    .A3(_03913_),
    .ZN(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09559_ (.A1(\as2650.stack[13][15] ),
    .A2(_03848_),
    .B1(_03849_),
    .B2(\as2650.stack[12][15] ),
    .ZN(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09560_ (.A1(\as2650.stack[14][15] ),
    .A2(_03832_),
    .B1(_03837_),
    .B2(\as2650.stack[15][15] ),
    .ZN(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09561_ (.A1(_03847_),
    .A2(_03915_),
    .A3(_03916_),
    .ZN(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09562_ (.A1(_03826_),
    .A2(_03914_),
    .A3(_03917_),
    .ZN(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09563_ (.A1(_03826_),
    .A2(_03911_),
    .B(_03918_),
    .ZN(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09564_ (.I0(_03919_),
    .I1(_02466_),
    .S(_03821_),
    .Z(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09565_ (.A1(_02466_),
    .A2(_03881_),
    .B1(_03920_),
    .B2(_03869_),
    .ZN(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09566_ (.A1(_03877_),
    .A2(_03921_),
    .B(_03817_),
    .ZN(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09567_ (.A1(_03877_),
    .A2(_03904_),
    .B(_03922_),
    .ZN(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09568_ (.A1(\as2650.instruction_args_latch[15] ),
    .A2(_03776_),
    .B(_01450_),
    .ZN(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09569_ (.A1(_03923_),
    .A2(_03924_),
    .ZN(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09570_ (.I(_01247_),
    .Z(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09571_ (.A1(\as2650.last_addr[8] ),
    .A2(_03925_),
    .ZN(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09572_ (.A1(_01551_),
    .A2(_03926_),
    .B(_03604_),
    .ZN(_00430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09573_ (.A1(_01207_),
    .A2(_01541_),
    .ZN(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09574_ (.A1(\as2650.last_addr[9] ),
    .A2(_03925_),
    .ZN(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09575_ (.A1(_03366_),
    .A2(_03927_),
    .A3(_03928_),
    .ZN(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09576_ (.A1(\as2650.last_addr[10] ),
    .A2(_03925_),
    .ZN(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09577_ (.A1(_01584_),
    .A2(_03929_),
    .B(_03357_),
    .ZN(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09578_ (.A1(\as2650.last_addr[11] ),
    .A2(_03925_),
    .ZN(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09579_ (.A1(_03366_),
    .A2(_01597_),
    .A3(_03930_),
    .ZN(_00433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09580_ (.A1(\as2650.last_addr[12] ),
    .A2(_01631_),
    .ZN(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09581_ (.A1(_01610_),
    .A2(_03931_),
    .B(_03357_),
    .ZN(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09582_ (.I(\as2650.last_addr[13] ),
    .ZN(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09583_ (.A1(_03932_),
    .A2(net204),
    .B(_03366_),
    .C(_01626_),
    .ZN(_00435_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09584_ (.A1(_01239_),
    .A2(_01631_),
    .Z(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09585_ (.A1(\as2650.last_addr[14] ),
    .A2(_01631_),
    .ZN(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09586_ (.A1(_03933_),
    .A2(_03934_),
    .B(_03357_),
    .ZN(_00436_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09587_ (.I(\as2650.last_addr[15] ),
    .ZN(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09588_ (.A1(_03935_),
    .A2(net204),
    .B(_03588_),
    .C(_01648_),
    .ZN(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09589_ (.I(_03621_),
    .Z(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09590_ (.I(_00912_),
    .Z(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _09591_ (.A1(_01504_),
    .A2(_02821_),
    .A3(_03937_),
    .A4(_01511_),
    .ZN(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09592_ (.A1(_03936_),
    .A2(_03938_),
    .ZN(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09593_ (.I(_03939_),
    .Z(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09594_ (.I(_03940_),
    .Z(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09595_ (.I(_03940_),
    .Z(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09596_ (.A1(\as2650.ivectors_base[0] ),
    .A2(_03942_),
    .ZN(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09597_ (.I(_01683_),
    .Z(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09598_ (.I(_03944_),
    .Z(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09599_ (.A1(_02317_),
    .A2(_03941_),
    .B(_03943_),
    .C(_03945_),
    .ZN(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09600_ (.A1(\as2650.ivectors_base[1] ),
    .A2(_03942_),
    .ZN(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09601_ (.A1(_02331_),
    .A2(_03941_),
    .B(_03946_),
    .C(_03945_),
    .ZN(_00439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09602_ (.A1(\as2650.ivectors_base[2] ),
    .A2(_03942_),
    .ZN(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09603_ (.A1(_02346_),
    .A2(_03941_),
    .B(_03947_),
    .C(_03945_),
    .ZN(_00440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09604_ (.A1(\as2650.ivectors_base[3] ),
    .A2(_03942_),
    .ZN(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09605_ (.A1(_02360_),
    .A2(_03941_),
    .B(_03948_),
    .C(_03945_),
    .ZN(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09606_ (.I(_03940_),
    .Z(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09607_ (.I(_03939_),
    .Z(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09608_ (.A1(\as2650.ivectors_base[4] ),
    .A2(_03950_),
    .ZN(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09609_ (.I(_03944_),
    .Z(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09610_ (.A1(_02376_),
    .A2(_03949_),
    .B(_03951_),
    .C(_03952_),
    .ZN(_00442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09611_ (.A1(\as2650.ivectors_base[5] ),
    .A2(_03950_),
    .ZN(_03953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09612_ (.A1(_02393_),
    .A2(_03949_),
    .B(_03953_),
    .C(_03952_),
    .ZN(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09613_ (.A1(\as2650.ivectors_base[6] ),
    .A2(_03950_),
    .ZN(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09614_ (.A1(_02406_),
    .A2(_03949_),
    .B(_03954_),
    .C(_03952_),
    .ZN(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09615_ (.A1(\as2650.ivectors_base[7] ),
    .A2(_03950_),
    .ZN(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09616_ (.A1(_02427_),
    .A2(_03949_),
    .B(_03955_),
    .C(_03952_),
    .ZN(_00445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09617_ (.I(_03940_),
    .Z(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09618_ (.I(_03939_),
    .Z(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09619_ (.A1(\as2650.ivectors_base[8] ),
    .A2(_03957_),
    .ZN(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09620_ (.I(_03944_),
    .Z(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09621_ (.A1(_02434_),
    .A2(_03956_),
    .B(_03958_),
    .C(_03959_),
    .ZN(_00446_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09622_ (.A1(\as2650.ivectors_base[9] ),
    .A2(_03957_),
    .ZN(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09623_ (.A1(_02451_),
    .A2(_03956_),
    .B(_03960_),
    .C(_03959_),
    .ZN(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09624_ (.A1(\as2650.ivectors_base[10] ),
    .A2(_03957_),
    .ZN(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09625_ (.A1(_02460_),
    .A2(_03956_),
    .B(_03961_),
    .C(_03959_),
    .ZN(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09626_ (.A1(\as2650.ivectors_base[11] ),
    .A2(_03957_),
    .ZN(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09627_ (.A1(_02469_),
    .A2(_03956_),
    .B(_03962_),
    .C(_03959_),
    .ZN(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09628_ (.I(_03716_),
    .Z(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09629_ (.I(_00947_),
    .Z(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09630_ (.I(_03964_),
    .Z(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09631_ (.A1(_02222_),
    .A2(_03965_),
    .ZN(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09632_ (.I(_03812_),
    .Z(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09633_ (.A1(_03966_),
    .A2(_03967_),
    .B(_03652_),
    .ZN(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _09634_ (.A1(_00660_),
    .A2(_02875_),
    .Z(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09635_ (.I(_01520_),
    .Z(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09636_ (.I(_03639_),
    .Z(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09637_ (.I(_03971_),
    .Z(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09638_ (.I(_02830_),
    .Z(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09639_ (.A1(_01659_),
    .A2(_03973_),
    .ZN(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09640_ (.A1(_02281_),
    .A2(_03974_),
    .Z(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09641_ (.I(_03819_),
    .Z(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09642_ (.I(_03822_),
    .Z(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09643_ (.A1(\as2650.stack[10][0] ),
    .A2(_02251_),
    .B1(_03834_),
    .B2(\as2650.stack[11][0] ),
    .ZN(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09644_ (.I(_02477_),
    .Z(_03979_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09645_ (.I(_02594_),
    .Z(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09646_ (.A1(\as2650.stack[9][0] ),
    .A2(_03979_),
    .B1(_03980_),
    .B2(\as2650.stack[8][0] ),
    .ZN(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09647_ (.A1(_03829_),
    .A2(_03978_),
    .A3(_03981_),
    .ZN(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09648_ (.I(_03843_),
    .Z(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09649_ (.A1(\as2650.stack[13][0] ),
    .A2(_03979_),
    .B1(_03980_),
    .B2(\as2650.stack[12][0] ),
    .ZN(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09650_ (.A1(\as2650.stack[14][0] ),
    .A2(_02251_),
    .B1(_03834_),
    .B2(\as2650.stack[15][0] ),
    .ZN(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09651_ (.A1(_03983_),
    .A2(_03984_),
    .A3(_03985_),
    .ZN(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09652_ (.A1(_03982_),
    .A2(_03986_),
    .Z(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09653_ (.I(_03844_),
    .Z(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09654_ (.I(_02250_),
    .Z(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09655_ (.I(_03833_),
    .Z(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09656_ (.I(_02476_),
    .Z(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09657_ (.I(_02593_),
    .Z(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09658_ (.A1(\as2650.stack[5][0] ),
    .A2(_03991_),
    .B1(_03992_),
    .B2(\as2650.stack[4][0] ),
    .ZN(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09659_ (.I(_03993_),
    .ZN(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09660_ (.A1(\as2650.stack[6][0] ),
    .A2(_03989_),
    .B1(_03990_),
    .B2(\as2650.stack[7][0] ),
    .C(_03994_),
    .ZN(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09661_ (.A1(_03988_),
    .A2(_03995_),
    .B(_03823_),
    .ZN(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09662_ (.I(_03828_),
    .Z(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09663_ (.I(_03997_),
    .Z(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09664_ (.I(_02249_),
    .Z(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09665_ (.I(_03999_),
    .Z(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09666_ (.I(_03827_),
    .Z(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09667_ (.I(_04001_),
    .Z(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09668_ (.A1(\as2650.stack[2][0] ),
    .A2(_04000_),
    .B1(_04002_),
    .B2(\as2650.stack[3][0] ),
    .ZN(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09669_ (.I(_02477_),
    .Z(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09670_ (.I(_04004_),
    .Z(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09671_ (.I(_02594_),
    .Z(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09672_ (.I(_04006_),
    .Z(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09673_ (.A1(\as2650.stack[1][0] ),
    .A2(_04005_),
    .B1(_04007_),
    .B2(\as2650.stack[0][0] ),
    .ZN(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09674_ (.A1(_03998_),
    .A2(_04003_),
    .A3(_04008_),
    .ZN(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _09675_ (.A1(_03977_),
    .A2(_03987_),
    .B1(_03996_),
    .B2(_04009_),
    .ZN(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09676_ (.A1(_03819_),
    .A2(_04010_),
    .ZN(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09677_ (.A1(_02281_),
    .A2(_03976_),
    .B(_04011_),
    .C(_03971_),
    .ZN(_04012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09678_ (.I(_01515_),
    .Z(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09679_ (.A1(_03972_),
    .A2(_03975_),
    .B(_04012_),
    .C(_04013_),
    .ZN(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09680_ (.A1(_02222_),
    .A2(_03970_),
    .B(_04014_),
    .ZN(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09681_ (.A1(_01680_),
    .A2(_04015_),
    .ZN(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09682_ (.I(_02863_),
    .Z(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09683_ (.I(_03413_),
    .Z(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09684_ (.A1(_03751_),
    .A2(_03414_),
    .ZN(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09685_ (.A1(_04018_),
    .A2(_03386_),
    .B(_03868_),
    .C(_04019_),
    .ZN(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09686_ (.I(_01225_),
    .Z(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09687_ (.A1(_04021_),
    .A2(_04015_),
    .ZN(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09688_ (.A1(_03615_),
    .A2(_03811_),
    .ZN(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09689_ (.I(_04023_),
    .Z(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09690_ (.A1(_03966_),
    .A2(_04022_),
    .B(_04024_),
    .ZN(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09691_ (.A1(_04017_),
    .A2(_04020_),
    .A3(_04025_),
    .ZN(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09692_ (.A1(_03969_),
    .A2(_04016_),
    .A3(_04026_),
    .ZN(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09693_ (.A1(_03400_),
    .A2(_03792_),
    .Z(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09694_ (.A1(_03968_),
    .A2(_04027_),
    .B1(_04028_),
    .B2(_03879_),
    .ZN(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09695_ (.A1(_03963_),
    .A2(_04029_),
    .ZN(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09696_ (.I(_03944_),
    .Z(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09697_ (.A1(_03752_),
    .A2(_03875_),
    .B(_04030_),
    .C(_04031_),
    .ZN(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09698_ (.A1(_03422_),
    .A2(_03790_),
    .Z(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09699_ (.A1(_04032_),
    .A2(_03793_),
    .Z(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09700_ (.A1(_03964_),
    .A2(_02283_),
    .ZN(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09701_ (.A1(_03967_),
    .A2(_04034_),
    .B(_03652_),
    .ZN(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09702_ (.A1(_00951_),
    .A2(_01406_),
    .A3(_01658_),
    .ZN(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09703_ (.A1(_02276_),
    .A2(_04036_),
    .Z(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09704_ (.I0(_02283_),
    .I1(_04037_),
    .S(_03699_),
    .Z(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09705_ (.A1(_02198_),
    .A2(_03738_),
    .ZN(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09706_ (.I(_04039_),
    .Z(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09707_ (.I(_03977_),
    .Z(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09708_ (.I(_03997_),
    .Z(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09709_ (.I(_02250_),
    .Z(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09710_ (.I(_04043_),
    .Z(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09711_ (.I(_03833_),
    .Z(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09712_ (.I(_04045_),
    .Z(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09713_ (.A1(\as2650.stack[2][1] ),
    .A2(_04044_),
    .B1(_04046_),
    .B2(\as2650.stack[3][1] ),
    .ZN(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09714_ (.I(_02478_),
    .Z(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09715_ (.I(_02595_),
    .Z(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09716_ (.A1(\as2650.stack[1][1] ),
    .A2(_04048_),
    .B1(_04049_),
    .B2(\as2650.stack[0][1] ),
    .ZN(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09717_ (.A1(_04042_),
    .A2(_04047_),
    .A3(_04050_),
    .ZN(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09718_ (.I(_03983_),
    .Z(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09719_ (.I(_02478_),
    .Z(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09720_ (.I(_02595_),
    .Z(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09721_ (.A1(\as2650.stack[5][1] ),
    .A2(_04053_),
    .B1(_04054_),
    .B2(\as2650.stack[4][1] ),
    .ZN(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09722_ (.I(_04043_),
    .Z(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09723_ (.I(_04045_),
    .Z(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09724_ (.A1(\as2650.stack[6][1] ),
    .A2(_04056_),
    .B1(_04057_),
    .B2(\as2650.stack[7][1] ),
    .ZN(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09725_ (.A1(_04052_),
    .A2(_04055_),
    .A3(_04058_),
    .ZN(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09726_ (.A1(_04051_),
    .A2(_04059_),
    .ZN(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09727_ (.I(_03823_),
    .Z(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09728_ (.I(_04043_),
    .Z(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09729_ (.I(_04045_),
    .Z(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09730_ (.A1(\as2650.stack[10][1] ),
    .A2(_04062_),
    .B1(_04063_),
    .B2(\as2650.stack[11][1] ),
    .ZN(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09731_ (.I(_04004_),
    .Z(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09732_ (.I(_04006_),
    .Z(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09733_ (.A1(\as2650.stack[9][1] ),
    .A2(_04065_),
    .B1(_04066_),
    .B2(\as2650.stack[8][1] ),
    .ZN(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09734_ (.A1(_04042_),
    .A2(_04064_),
    .A3(_04067_),
    .ZN(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09735_ (.A1(\as2650.stack[13][1] ),
    .A2(_04065_),
    .B1(_04066_),
    .B2(\as2650.stack[12][1] ),
    .ZN(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09736_ (.A1(\as2650.stack[14][1] ),
    .A2(_04062_),
    .B1(_04063_),
    .B2(\as2650.stack[15][1] ),
    .ZN(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09737_ (.A1(_03845_),
    .A2(_04069_),
    .A3(_04070_),
    .ZN(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09738_ (.A1(_04061_),
    .A2(_04068_),
    .A3(_04071_),
    .ZN(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09739_ (.A1(_04041_),
    .A2(_04060_),
    .B(_04072_),
    .ZN(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09740_ (.I(_04039_),
    .Z(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09741_ (.A1(_02283_),
    .A2(_04074_),
    .ZN(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09742_ (.A1(_04040_),
    .A2(_04073_),
    .B(_04075_),
    .C(_03640_),
    .ZN(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09743_ (.A1(_03972_),
    .A2(_04038_),
    .B(_04076_),
    .C(_04013_),
    .ZN(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09744_ (.A1(_02276_),
    .A2(_03970_),
    .B(_04077_),
    .ZN(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09745_ (.A1(_01680_),
    .A2(_04078_),
    .ZN(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09746_ (.I(_03867_),
    .Z(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09747_ (.A1(_04021_),
    .A2(_04078_),
    .ZN(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09748_ (.A1(_04034_),
    .A2(_04081_),
    .ZN(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09749_ (.A1(_03416_),
    .A2(_04080_),
    .ZN(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09750_ (.A1(_04080_),
    .A2(_04082_),
    .B(_04083_),
    .C(_04017_),
    .ZN(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09751_ (.A1(_03969_),
    .A2(_04079_),
    .A3(_04084_),
    .ZN(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09752_ (.A1(_03879_),
    .A2(_04033_),
    .B1(_04035_),
    .B2(_04085_),
    .ZN(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09753_ (.A1(_03963_),
    .A2(_04086_),
    .ZN(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09754_ (.A1(_03757_),
    .A2(_03875_),
    .B(_04087_),
    .C(_04031_),
    .ZN(_00451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09755_ (.I(_03747_),
    .Z(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09756_ (.I(_03818_),
    .Z(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09757_ (.A1(net189),
    .A2(_03806_),
    .ZN(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09758_ (.A1(_03437_),
    .A2(_04090_),
    .Z(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09759_ (.A1(_03795_),
    .A2(_04091_),
    .Z(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09760_ (.I(_03721_),
    .Z(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09761_ (.I(_01225_),
    .Z(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09762_ (.I(_04094_),
    .Z(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09763_ (.I(_03812_),
    .Z(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09764_ (.I(_04096_),
    .Z(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09765_ (.A1(_04095_),
    .A2(_03448_),
    .B(_04097_),
    .ZN(_04098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09766_ (.I(_03679_),
    .Z(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09767_ (.I(_04074_),
    .Z(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09768_ (.I(_03977_),
    .Z(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09769_ (.I(_03989_),
    .Z(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09770_ (.I(_03990_),
    .Z(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09771_ (.A1(\as2650.stack[10][2] ),
    .A2(_04102_),
    .B1(_04103_),
    .B2(\as2650.stack[11][2] ),
    .ZN(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09772_ (.I(_03979_),
    .Z(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09773_ (.I(_03980_),
    .Z(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09774_ (.A1(\as2650.stack[9][2] ),
    .A2(_04105_),
    .B1(_04106_),
    .B2(\as2650.stack[8][2] ),
    .ZN(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09775_ (.A1(_03830_),
    .A2(_04104_),
    .A3(_04107_),
    .ZN(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09776_ (.I(_03983_),
    .Z(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09777_ (.A1(\as2650.stack[13][2] ),
    .A2(_04105_),
    .B1(_04106_),
    .B2(\as2650.stack[12][2] ),
    .ZN(_04110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09778_ (.A1(\as2650.stack[14][2] ),
    .A2(_04102_),
    .B1(_04103_),
    .B2(\as2650.stack[15][2] ),
    .ZN(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09779_ (.A1(_04109_),
    .A2(_04110_),
    .A3(_04111_),
    .ZN(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09780_ (.A1(_04108_),
    .A2(_04112_),
    .Z(_04113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09781_ (.I(_03988_),
    .Z(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09782_ (.I(_02250_),
    .Z(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09783_ (.I(_04115_),
    .Z(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09784_ (.I(_03833_),
    .Z(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09785_ (.I(_04117_),
    .Z(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09786_ (.I(_03991_),
    .Z(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09787_ (.I(_03992_),
    .Z(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09788_ (.A1(\as2650.stack[5][2] ),
    .A2(_04119_),
    .B1(_04120_),
    .B2(\as2650.stack[4][2] ),
    .ZN(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09789_ (.I(_04121_),
    .ZN(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09790_ (.A1(\as2650.stack[6][2] ),
    .A2(_04116_),
    .B1(_04118_),
    .B2(\as2650.stack[7][2] ),
    .C(_04122_),
    .ZN(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09791_ (.A1(_04114_),
    .A2(_04123_),
    .B(_04041_),
    .ZN(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09792_ (.I(_03998_),
    .Z(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09793_ (.I(_04115_),
    .Z(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09794_ (.I(_04117_),
    .Z(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09795_ (.A1(\as2650.stack[2][2] ),
    .A2(_04126_),
    .B1(_04127_),
    .B2(\as2650.stack[3][2] ),
    .ZN(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09796_ (.I(_04119_),
    .Z(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09797_ (.I(_04120_),
    .Z(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09798_ (.A1(\as2650.stack[1][2] ),
    .A2(_04129_),
    .B1(_04130_),
    .B2(\as2650.stack[0][2] ),
    .ZN(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09799_ (.A1(_04125_),
    .A2(_04128_),
    .A3(_04131_),
    .ZN(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _09800_ (.A1(_04101_),
    .A2(_04113_),
    .B1(_04124_),
    .B2(_04132_),
    .ZN(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09801_ (.I(_04074_),
    .Z(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09802_ (.A1(_03448_),
    .A2(_04134_),
    .ZN(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09803_ (.A1(_04100_),
    .A2(_04133_),
    .B(_04135_),
    .C(_03972_),
    .ZN(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09804_ (.I(_03699_),
    .Z(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09805_ (.I(_03973_),
    .Z(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09806_ (.A1(_02275_),
    .A2(_04036_),
    .Z(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09807_ (.A1(_02296_),
    .A2(_04139_),
    .Z(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09808_ (.A1(_04138_),
    .A2(_04140_),
    .B(_03640_),
    .ZN(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09809_ (.A1(_02298_),
    .A2(_04137_),
    .B(_04141_),
    .ZN(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09810_ (.A1(_03629_),
    .A2(_04136_),
    .A3(_04142_),
    .ZN(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09811_ (.A1(_02296_),
    .A2(_03936_),
    .ZN(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09812_ (.A1(_04143_),
    .A2(_04144_),
    .ZN(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09813_ (.I(_03969_),
    .Z(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09814_ (.A1(_04099_),
    .A2(_04145_),
    .B(_04146_),
    .ZN(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09815_ (.I(_03868_),
    .Z(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09816_ (.I(_01225_),
    .Z(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09817_ (.A1(_04149_),
    .A2(_03448_),
    .ZN(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09818_ (.I(_00947_),
    .Z(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09819_ (.A1(_04151_),
    .A2(_04145_),
    .ZN(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09820_ (.A1(_04150_),
    .A2(_04152_),
    .B(_04080_),
    .ZN(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09821_ (.I(_03722_),
    .Z(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09822_ (.A1(_03434_),
    .A2(_04148_),
    .B(_04153_),
    .C(_04154_),
    .ZN(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09823_ (.A1(_04093_),
    .A2(_04098_),
    .B1(_04147_),
    .B2(_04155_),
    .ZN(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09824_ (.A1(_04089_),
    .A2(_04092_),
    .B(_04156_),
    .ZN(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09825_ (.I(_03746_),
    .Z(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09826_ (.I(_01449_),
    .Z(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09827_ (.A1(_03660_),
    .A2(_04158_),
    .B(_04159_),
    .ZN(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09828_ (.A1(_04088_),
    .A2(_04157_),
    .B(_04160_),
    .ZN(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09829_ (.I(_03717_),
    .Z(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09830_ (.I(_04017_),
    .Z(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09831_ (.I(_04024_),
    .Z(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09832_ (.I(_04021_),
    .Z(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09833_ (.I(_04013_),
    .Z(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09834_ (.I(_03640_),
    .Z(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09835_ (.A1(_02311_),
    .A2(_04137_),
    .ZN(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09836_ (.I(_03973_),
    .ZN(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09837_ (.I(_04168_),
    .Z(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09838_ (.A1(_02295_),
    .A2(\as2650.PC[3] ),
    .A3(_04139_),
    .Z(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09839_ (.A1(_02296_),
    .A2(_04139_),
    .B(_02306_),
    .ZN(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09840_ (.A1(_04169_),
    .A2(_04170_),
    .A3(_04171_),
    .ZN(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09841_ (.I(_03819_),
    .Z(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09842_ (.A1(\as2650.stack[2][3] ),
    .A2(_04056_),
    .B1(_04057_),
    .B2(\as2650.stack[3][3] ),
    .ZN(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09843_ (.A1(\as2650.stack[1][3] ),
    .A2(_04048_),
    .B1(_04049_),
    .B2(\as2650.stack[0][3] ),
    .ZN(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09844_ (.A1(_04042_),
    .A2(_04174_),
    .A3(_04175_),
    .ZN(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09845_ (.A1(\as2650.stack[5][3] ),
    .A2(_04053_),
    .B1(_04054_),
    .B2(\as2650.stack[4][3] ),
    .ZN(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09846_ (.A1(\as2650.stack[6][3] ),
    .A2(_04056_),
    .B1(_04057_),
    .B2(\as2650.stack[7][3] ),
    .ZN(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09847_ (.A1(_04052_),
    .A2(_04177_),
    .A3(_04178_),
    .ZN(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09848_ (.A1(_04176_),
    .A2(_04179_),
    .ZN(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09849_ (.A1(\as2650.stack[10][3] ),
    .A2(_04000_),
    .B1(_04063_),
    .B2(\as2650.stack[11][3] ),
    .ZN(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09850_ (.A1(\as2650.stack[9][3] ),
    .A2(_04065_),
    .B1(_04066_),
    .B2(\as2650.stack[8][3] ),
    .ZN(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09851_ (.A1(_03998_),
    .A2(_04181_),
    .A3(_04182_),
    .ZN(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09852_ (.A1(\as2650.stack[13][3] ),
    .A2(_04065_),
    .B1(_04066_),
    .B2(\as2650.stack[12][3] ),
    .ZN(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09853_ (.A1(\as2650.stack[14][3] ),
    .A2(_04062_),
    .B1(_04002_),
    .B2(\as2650.stack[15][3] ),
    .ZN(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09854_ (.A1(_03845_),
    .A2(_04184_),
    .A3(_04185_),
    .ZN(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09855_ (.A1(_04061_),
    .A2(_04183_),
    .A3(_04186_),
    .ZN(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09856_ (.A1(_04041_),
    .A2(_04180_),
    .B(_04187_),
    .ZN(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09857_ (.A1(_03976_),
    .A2(_04188_),
    .ZN(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09858_ (.I(_03639_),
    .Z(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09859_ (.A1(_02311_),
    .A2(_04173_),
    .B(_04189_),
    .C(_04190_),
    .ZN(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09860_ (.A1(_04166_),
    .A2(_04167_),
    .A3(_04172_),
    .B(_04191_),
    .ZN(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09861_ (.A1(_04165_),
    .A2(_04192_),
    .ZN(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09862_ (.A1(_02306_),
    .A2(_03630_),
    .B(_04193_),
    .ZN(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09863_ (.A1(_03965_),
    .A2(_02311_),
    .Z(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09864_ (.I(_04023_),
    .Z(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09865_ (.A1(_04164_),
    .A2(_04194_),
    .B(_04195_),
    .C(_04196_),
    .ZN(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09866_ (.A1(_03457_),
    .A2(_04163_),
    .B(_04197_),
    .ZN(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09867_ (.A1(_04162_),
    .A2(_04198_),
    .ZN(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09868_ (.A1(_04149_),
    .A2(_04096_),
    .B(_03392_),
    .ZN(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09869_ (.A1(_01681_),
    .A2(_04194_),
    .ZN(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09870_ (.A1(_04199_),
    .A2(_04200_),
    .A3(_04201_),
    .ZN(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09871_ (.A1(_03721_),
    .A2(_04096_),
    .Z(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09872_ (.A1(_04195_),
    .A2(_04203_),
    .B(_03899_),
    .ZN(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09873_ (.A1(_03788_),
    .A2(_03797_),
    .B(_03814_),
    .ZN(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09874_ (.A1(_03788_),
    .A2(_03797_),
    .B(_04205_),
    .ZN(_04206_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09875_ (.A1(_04204_),
    .A2(_04206_),
    .ZN(_04207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09876_ (.A1(_03762_),
    .A2(_04161_),
    .B1(_04202_),
    .B2(_04207_),
    .C(_03517_),
    .ZN(_00453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09877_ (.A1(net191),
    .A2(_03806_),
    .ZN(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09878_ (.A1(_03482_),
    .A2(_04208_),
    .Z(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09879_ (.A1(_03799_),
    .A2(_04209_),
    .Z(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09880_ (.A1(_04095_),
    .A2(_03489_),
    .B(_04097_),
    .ZN(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09881_ (.I(_03829_),
    .Z(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09882_ (.A1(\as2650.stack[2][4] ),
    .A2(_04116_),
    .B1(_04118_),
    .B2(\as2650.stack[3][4] ),
    .ZN(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09883_ (.I(_04119_),
    .Z(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09884_ (.I(_04120_),
    .Z(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09885_ (.A1(\as2650.stack[1][4] ),
    .A2(_04214_),
    .B1(_04215_),
    .B2(\as2650.stack[0][4] ),
    .ZN(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09886_ (.A1(_04212_),
    .A2(_04213_),
    .A3(_04216_),
    .ZN(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09887_ (.A1(\as2650.stack[5][4] ),
    .A2(_04214_),
    .B1(_04215_),
    .B2(\as2650.stack[4][4] ),
    .ZN(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09888_ (.I(_04115_),
    .Z(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09889_ (.I(_04117_),
    .Z(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09890_ (.A1(\as2650.stack[6][4] ),
    .A2(_04219_),
    .B1(_04220_),
    .B2(\as2650.stack[7][4] ),
    .ZN(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09891_ (.A1(_04114_),
    .A2(_04218_),
    .A3(_04221_),
    .ZN(_04222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09892_ (.A1(_04217_),
    .A2(_04222_),
    .ZN(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09893_ (.A1(\as2650.stack[10][4] ),
    .A2(_04116_),
    .B1(_04118_),
    .B2(\as2650.stack[11][4] ),
    .ZN(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09894_ (.A1(\as2650.stack[9][4] ),
    .A2(_04214_),
    .B1(_04215_),
    .B2(\as2650.stack[8][4] ),
    .ZN(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09895_ (.A1(_04212_),
    .A2(_04224_),
    .A3(_04225_),
    .ZN(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09896_ (.A1(\as2650.stack[13][4] ),
    .A2(_04214_),
    .B1(_04215_),
    .B2(\as2650.stack[12][4] ),
    .ZN(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09897_ (.A1(\as2650.stack[14][4] ),
    .A2(_04219_),
    .B1(_04220_),
    .B2(\as2650.stack[15][4] ),
    .ZN(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09898_ (.A1(_04114_),
    .A2(_04227_),
    .A3(_04228_),
    .ZN(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09899_ (.A1(_04226_),
    .A2(_04229_),
    .ZN(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _09900_ (.I0(_04223_),
    .I1(_04230_),
    .S(_03824_),
    .Z(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09901_ (.A1(_03489_),
    .A2(_04134_),
    .ZN(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09902_ (.I(_03971_),
    .Z(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09903_ (.A1(_04100_),
    .A2(_04231_),
    .B(_04232_),
    .C(_04233_),
    .ZN(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09904_ (.A1(_02322_),
    .A2(_04170_),
    .Z(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09905_ (.I(_03639_),
    .Z(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09906_ (.A1(_04138_),
    .A2(_04235_),
    .B(_04236_),
    .ZN(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09907_ (.A1(_02324_),
    .A2(_03700_),
    .B(_04237_),
    .ZN(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09908_ (.A1(_04234_),
    .A2(_04238_),
    .ZN(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09909_ (.A1(_02322_),
    .A2(_03936_),
    .ZN(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09910_ (.A1(_03622_),
    .A2(_04239_),
    .B(_04240_),
    .ZN(_04241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09911_ (.A1(_04099_),
    .A2(_04241_),
    .B(_04146_),
    .ZN(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09912_ (.I0(_03489_),
    .I1(_04241_),
    .S(_03965_),
    .Z(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09913_ (.I(_04023_),
    .Z(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09914_ (.A1(_03455_),
    .A2(_03478_),
    .ZN(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09915_ (.A1(_03182_),
    .A2(_03454_),
    .B(_04244_),
    .C(_04245_),
    .ZN(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09916_ (.I(_01679_),
    .Z(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09917_ (.A1(_04163_),
    .A2(_04243_),
    .B(_04246_),
    .C(_04247_),
    .ZN(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09918_ (.A1(_04093_),
    .A2(_04211_),
    .B1(_04242_),
    .B2(_04248_),
    .ZN(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09919_ (.A1(_04089_),
    .A2(_04210_),
    .B(_04249_),
    .ZN(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09920_ (.A1(_03663_),
    .A2(_04158_),
    .B(_04159_),
    .ZN(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09921_ (.A1(_04088_),
    .A2(_04250_),
    .B(_04251_),
    .ZN(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09922_ (.A1(_02338_),
    .A2(_04137_),
    .ZN(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09923_ (.I(_04168_),
    .Z(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _09924_ (.A1(_02321_),
    .A2(_02334_),
    .A3(_04170_),
    .Z(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09925_ (.A1(_02322_),
    .A2(_04170_),
    .B(_02335_),
    .ZN(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09926_ (.A1(_04253_),
    .A2(_04254_),
    .A3(_04255_),
    .ZN(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09927_ (.I(_03822_),
    .Z(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09928_ (.A1(\as2650.stack[2][5] ),
    .A2(_04056_),
    .B1(_04057_),
    .B2(\as2650.stack[3][5] ),
    .ZN(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09929_ (.A1(\as2650.stack[1][5] ),
    .A2(_04053_),
    .B1(_04054_),
    .B2(\as2650.stack[0][5] ),
    .ZN(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09930_ (.A1(_04042_),
    .A2(_04258_),
    .A3(_04259_),
    .ZN(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09931_ (.A1(\as2650.stack[5][5] ),
    .A2(_04053_),
    .B1(_04054_),
    .B2(\as2650.stack[4][5] ),
    .ZN(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09932_ (.A1(\as2650.stack[6][5] ),
    .A2(_04062_),
    .B1(_04063_),
    .B2(\as2650.stack[7][5] ),
    .ZN(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09933_ (.A1(_03845_),
    .A2(_04261_),
    .A3(_04262_),
    .ZN(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09934_ (.A1(_04260_),
    .A2(_04263_),
    .ZN(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09935_ (.A1(\as2650.stack[10][5] ),
    .A2(_04000_),
    .B1(_04002_),
    .B2(\as2650.stack[11][5] ),
    .ZN(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09936_ (.A1(\as2650.stack[9][5] ),
    .A2(_04005_),
    .B1(_04007_),
    .B2(\as2650.stack[8][5] ),
    .ZN(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09937_ (.A1(_03998_),
    .A2(_04265_),
    .A3(_04266_),
    .ZN(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09938_ (.A1(\as2650.stack[13][5] ),
    .A2(_04005_),
    .B1(_04007_),
    .B2(\as2650.stack[12][5] ),
    .ZN(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09939_ (.A1(\as2650.stack[14][5] ),
    .A2(_04000_),
    .B1(_04002_),
    .B2(\as2650.stack[15][5] ),
    .ZN(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09940_ (.A1(_03988_),
    .A2(_04268_),
    .A3(_04269_),
    .ZN(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09941_ (.A1(_04061_),
    .A2(_04267_),
    .A3(_04270_),
    .ZN(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09942_ (.A1(_04257_),
    .A2(_04264_),
    .B(_04271_),
    .ZN(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09943_ (.A1(_03976_),
    .A2(_04272_),
    .ZN(_04273_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09944_ (.A1(_02338_),
    .A2(_04173_),
    .B(_04273_),
    .C(_04190_),
    .ZN(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09945_ (.A1(_04166_),
    .A2(_04252_),
    .A3(_04256_),
    .B(_04274_),
    .ZN(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09946_ (.A1(_04165_),
    .A2(_04275_),
    .ZN(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09947_ (.A1(_02335_),
    .A2(_03630_),
    .B(_04276_),
    .ZN(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09948_ (.A1(_04094_),
    .A2(_03485_),
    .ZN(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09949_ (.A1(_04164_),
    .A2(_04277_),
    .B(_04278_),
    .C(_04196_),
    .ZN(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09950_ (.A1(_03495_),
    .A2(_04163_),
    .B(_04279_),
    .ZN(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09951_ (.A1(_04162_),
    .A2(_04280_),
    .ZN(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09952_ (.I(_03722_),
    .Z(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09953_ (.A1(_04282_),
    .A2(_04277_),
    .ZN(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09954_ (.A1(_04200_),
    .A2(_04281_),
    .A3(_04283_),
    .ZN(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09955_ (.A1(_03785_),
    .A2(_03801_),
    .B(_03876_),
    .ZN(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09956_ (.A1(_03785_),
    .A2(_03801_),
    .B(_04285_),
    .ZN(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09957_ (.A1(_04203_),
    .A2(_04278_),
    .B(_03899_),
    .ZN(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09958_ (.A1(_04286_),
    .A2(_04287_),
    .ZN(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09959_ (.A1(_03768_),
    .A2(_04161_),
    .B1(_04284_),
    .B2(_04288_),
    .C(_01446_),
    .ZN(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09960_ (.I(_01520_),
    .Z(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09961_ (.A1(\as2650.stack[2][6] ),
    .A2(_04043_),
    .B1(_04045_),
    .B2(\as2650.stack[3][6] ),
    .ZN(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09962_ (.A1(\as2650.stack[1][6] ),
    .A2(_04004_),
    .B1(_04006_),
    .B2(\as2650.stack[0][6] ),
    .ZN(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09963_ (.A1(_03997_),
    .A2(_04290_),
    .A3(_04291_),
    .ZN(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09964_ (.A1(\as2650.stack[5][6] ),
    .A2(_04004_),
    .B1(_04006_),
    .B2(\as2650.stack[4][6] ),
    .ZN(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09965_ (.A1(\as2650.stack[6][6] ),
    .A2(_03999_),
    .B1(_04001_),
    .B2(\as2650.stack[7][6] ),
    .ZN(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09966_ (.A1(_03844_),
    .A2(_04293_),
    .A3(_04294_),
    .ZN(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09967_ (.A1(_04292_),
    .A2(_04295_),
    .ZN(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09968_ (.A1(\as2650.stack[10][6] ),
    .A2(_03999_),
    .B1(_04001_),
    .B2(\as2650.stack[11][6] ),
    .ZN(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09969_ (.A1(\as2650.stack[9][6] ),
    .A2(_03991_),
    .B1(_03992_),
    .B2(\as2650.stack[8][6] ),
    .ZN(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09970_ (.A1(_03828_),
    .A2(_04297_),
    .A3(_04298_),
    .ZN(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09971_ (.A1(\as2650.stack[13][6] ),
    .A2(_03991_),
    .B1(_03992_),
    .B2(\as2650.stack[12][6] ),
    .ZN(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09972_ (.A1(\as2650.stack[14][6] ),
    .A2(_03999_),
    .B1(_04001_),
    .B2(\as2650.stack[15][6] ),
    .ZN(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09973_ (.A1(_03844_),
    .A2(_04300_),
    .A3(_04301_),
    .ZN(_04302_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09974_ (.A1(_03822_),
    .A2(_04299_),
    .A3(_04302_),
    .ZN(_04303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09975_ (.A1(_03823_),
    .A2(_04296_),
    .B(_04303_),
    .ZN(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09976_ (.A1(_04134_),
    .A2(_04304_),
    .Z(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09977_ (.A1(_02354_),
    .A2(_03820_),
    .B(_04305_),
    .C(_04233_),
    .ZN(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09978_ (.A1(_02351_),
    .A2(_04254_),
    .ZN(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09979_ (.A1(_04137_),
    .A2(_04307_),
    .B(_04190_),
    .ZN(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09980_ (.A1(_02354_),
    .A2(_03700_),
    .B(_04308_),
    .ZN(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09981_ (.A1(_04289_),
    .A2(_04306_),
    .A3(_04309_),
    .ZN(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09982_ (.A1(_02351_),
    .A2(_03643_),
    .B(_04310_),
    .ZN(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09983_ (.A1(_04094_),
    .A2(_02354_),
    .ZN(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09984_ (.A1(_04164_),
    .A2(_04311_),
    .B(_04312_),
    .C(_04244_),
    .ZN(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09985_ (.A1(_03241_),
    .A2(_03414_),
    .ZN(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09986_ (.A1(_04018_),
    .A2(_03509_),
    .B(_04314_),
    .ZN(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09987_ (.A1(_04148_),
    .A2(_04315_),
    .ZN(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09988_ (.A1(_04313_),
    .A2(_04316_),
    .B(_04247_),
    .ZN(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09989_ (.I(_04200_),
    .ZN(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09990_ (.A1(_04282_),
    .A2(_04311_),
    .B(_04317_),
    .C(_04318_),
    .ZN(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09991_ (.A1(net194),
    .A2(_03806_),
    .ZN(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09992_ (.A1(_03514_),
    .A2(_04320_),
    .ZN(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09993_ (.A1(_03803_),
    .A2(_04321_),
    .Z(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09994_ (.A1(_04203_),
    .A2(_04312_),
    .B1(_04322_),
    .B2(_03818_),
    .C(_03899_),
    .ZN(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09995_ (.A1(_03672_),
    .A2(_03776_),
    .B1(_04319_),
    .B2(_04323_),
    .ZN(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09996_ (.A1(_03775_),
    .A2(_04324_),
    .ZN(_00456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09997_ (.A1(_02351_),
    .A2(_04254_),
    .ZN(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09998_ (.A1(_02364_),
    .A2(_04325_),
    .Z(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09999_ (.A1(_02368_),
    .A2(_04253_),
    .ZN(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10000_ (.A1(_04169_),
    .A2(_04326_),
    .B(_04327_),
    .ZN(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10001_ (.I(_04074_),
    .Z(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10002_ (.I(_03997_),
    .Z(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10003_ (.A1(\as2650.stack[10][7] ),
    .A2(_02252_),
    .B1(_03835_),
    .B2(\as2650.stack[11][7] ),
    .ZN(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10004_ (.A1(\as2650.stack[9][7] ),
    .A2(_02479_),
    .B1(_02596_),
    .B2(\as2650.stack[8][7] ),
    .ZN(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10005_ (.A1(_04330_),
    .A2(_04331_),
    .A3(_04332_),
    .ZN(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10006_ (.A1(\as2650.stack[13][7] ),
    .A2(_02479_),
    .B1(_02596_),
    .B2(\as2650.stack[12][7] ),
    .ZN(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10007_ (.A1(\as2650.stack[14][7] ),
    .A2(_02252_),
    .B1(_03835_),
    .B2(\as2650.stack[15][7] ),
    .ZN(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10008_ (.A1(_04052_),
    .A2(_04334_),
    .A3(_04335_),
    .ZN(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10009_ (.A1(_04333_),
    .A2(_04336_),
    .Z(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10010_ (.I(_03989_),
    .Z(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10011_ (.I(_03990_),
    .Z(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10012_ (.I(_02477_),
    .Z(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10013_ (.I(_02594_),
    .Z(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10014_ (.A1(\as2650.stack[5][7] ),
    .A2(_04340_),
    .B1(_04341_),
    .B2(\as2650.stack[4][7] ),
    .ZN(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10015_ (.I(_04342_),
    .ZN(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10016_ (.A1(\as2650.stack[6][7] ),
    .A2(_04338_),
    .B1(_04339_),
    .B2(\as2650.stack[7][7] ),
    .C(_04343_),
    .ZN(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10017_ (.A1(_04114_),
    .A2(_04344_),
    .B(_04257_),
    .ZN(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10018_ (.A1(\as2650.stack[2][7] ),
    .A2(_04126_),
    .B1(_04127_),
    .B2(\as2650.stack[3][7] ),
    .ZN(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10019_ (.A1(\as2650.stack[1][7] ),
    .A2(_04129_),
    .B1(_04130_),
    .B2(\as2650.stack[0][7] ),
    .ZN(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10020_ (.A1(_04125_),
    .A2(_04346_),
    .A3(_04347_),
    .ZN(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _10021_ (.A1(_04101_),
    .A2(_04337_),
    .B1(_04345_),
    .B2(_04348_),
    .ZN(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10022_ (.A1(_02368_),
    .A2(_04040_),
    .ZN(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10023_ (.A1(_04329_),
    .A2(_04349_),
    .B(_04350_),
    .C(_04236_),
    .ZN(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10024_ (.A1(_04166_),
    .A2(_04328_),
    .B(_04351_),
    .ZN(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10025_ (.A1(_04289_),
    .A2(_04352_),
    .ZN(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10026_ (.A1(_02364_),
    .A2(_03643_),
    .B(_04353_),
    .ZN(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10027_ (.A1(_04021_),
    .A2(_02368_),
    .ZN(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10028_ (.A1(_04149_),
    .A2(_04354_),
    .B(_04355_),
    .C(_04244_),
    .ZN(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10029_ (.A1(_04018_),
    .A2(_03524_),
    .B(_04314_),
    .ZN(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10030_ (.A1(_04080_),
    .A2(_04357_),
    .ZN(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10031_ (.A1(_04356_),
    .A2(_04358_),
    .B(_04247_),
    .ZN(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10032_ (.A1(_04282_),
    .A2(_04354_),
    .B(_04359_),
    .C(_04318_),
    .ZN(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10033_ (.A1(_04203_),
    .A2(_04355_),
    .B(_03817_),
    .ZN(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10034_ (.A1(_03781_),
    .A2(_03805_),
    .B(_03814_),
    .ZN(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10035_ (.A1(_03781_),
    .A2(_03805_),
    .B(_04362_),
    .ZN(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _10036_ (.A1(_04360_),
    .A2(_04361_),
    .A3(_04363_),
    .B1(_03747_),
    .B2(_03675_),
    .ZN(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10037_ (.A1(_03775_),
    .A2(_04364_),
    .ZN(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10038_ (.A1(_03777_),
    .A2(_03808_),
    .Z(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10039_ (.A1(_04095_),
    .A2(_02384_),
    .B(_03967_),
    .ZN(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10040_ (.A1(_04093_),
    .A2(_04366_),
    .ZN(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10041_ (.A1(_02350_),
    .A2(_02364_),
    .A3(_04254_),
    .ZN(_04368_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10042_ (.A1(_02385_),
    .A2(_04368_),
    .Z(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10043_ (.A1(_02384_),
    .A2(_04253_),
    .ZN(_04370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10044_ (.A1(_04169_),
    .A2(_04369_),
    .B(_04370_),
    .ZN(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10045_ (.A1(\as2650.stack[10][8] ),
    .A2(_04102_),
    .B1(_04103_),
    .B2(\as2650.stack[11][8] ),
    .ZN(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10046_ (.A1(\as2650.stack[9][8] ),
    .A2(_04105_),
    .B1(_04106_),
    .B2(\as2650.stack[8][8] ),
    .ZN(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10047_ (.A1(_03830_),
    .A2(_04372_),
    .A3(_04373_),
    .ZN(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10048_ (.I(_03983_),
    .Z(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10049_ (.A1(\as2650.stack[13][8] ),
    .A2(_04105_),
    .B1(_04106_),
    .B2(\as2650.stack[12][8] ),
    .ZN(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10050_ (.A1(\as2650.stack[14][8] ),
    .A2(_04102_),
    .B1(_04103_),
    .B2(\as2650.stack[15][8] ),
    .ZN(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10051_ (.A1(_04375_),
    .A2(_04376_),
    .A3(_04377_),
    .ZN(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10052_ (.A1(_04374_),
    .A2(_04378_),
    .Z(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10053_ (.A1(\as2650.stack[5][8] ),
    .A2(_04005_),
    .B1(_04007_),
    .B2(\as2650.stack[4][8] ),
    .ZN(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10054_ (.I(_04380_),
    .ZN(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10055_ (.A1(\as2650.stack[6][8] ),
    .A2(_04126_),
    .B1(_04127_),
    .B2(\as2650.stack[7][8] ),
    .C(_04381_),
    .ZN(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10056_ (.A1(_03846_),
    .A2(_04382_),
    .B(_04041_),
    .ZN(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10057_ (.A1(\as2650.stack[2][8] ),
    .A2(_04126_),
    .B1(_04127_),
    .B2(\as2650.stack[3][8] ),
    .ZN(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10058_ (.A1(\as2650.stack[1][8] ),
    .A2(_04129_),
    .B1(_04130_),
    .B2(\as2650.stack[0][8] ),
    .ZN(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10059_ (.A1(_04125_),
    .A2(_04384_),
    .A3(_04385_),
    .ZN(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _10060_ (.A1(_04101_),
    .A2(_04379_),
    .B1(_04383_),
    .B2(_04386_),
    .ZN(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10061_ (.A1(_02383_),
    .A2(_04040_),
    .ZN(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10062_ (.A1(_04329_),
    .A2(_04387_),
    .B(_04388_),
    .C(_04190_),
    .ZN(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10063_ (.A1(_03641_),
    .A2(_04371_),
    .B(_04389_),
    .ZN(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10064_ (.A1(_04165_),
    .A2(_04390_),
    .ZN(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10065_ (.A1(_02385_),
    .A2(_03643_),
    .B(_04391_),
    .ZN(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10066_ (.A1(_04094_),
    .A2(_02384_),
    .ZN(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10067_ (.A1(_04164_),
    .A2(_04392_),
    .B(_04393_),
    .C(_04244_),
    .ZN(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10068_ (.A1(_04018_),
    .A2(_03538_),
    .B(_04314_),
    .ZN(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10069_ (.A1(_04148_),
    .A2(_04395_),
    .ZN(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10070_ (.A1(_04394_),
    .A2(_04396_),
    .B(_04247_),
    .ZN(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10071_ (.A1(_00660_),
    .A2(_03721_),
    .ZN(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10072_ (.A1(_04282_),
    .A2(_04392_),
    .B(_04397_),
    .C(_04398_),
    .ZN(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10073_ (.A1(_04089_),
    .A2(_04365_),
    .B1(_04367_),
    .B2(_04399_),
    .ZN(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10074_ (.I(_01449_),
    .Z(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10075_ (.A1(\as2650.instruction_args_latch[8] ),
    .A2(_04158_),
    .B(_04401_),
    .ZN(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10076_ (.A1(_04088_),
    .A2(_04400_),
    .B(_04402_),
    .ZN(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10077_ (.A1(_03777_),
    .A2(_03808_),
    .Z(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10078_ (.A1(_03409_),
    .A2(_04403_),
    .ZN(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10079_ (.A1(_03409_),
    .A2(_04403_),
    .Z(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10080_ (.A1(_04404_),
    .A2(_04405_),
    .B(_03879_),
    .ZN(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10081_ (.A1(_04095_),
    .A2(_02399_),
    .B(_03967_),
    .ZN(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10082_ (.A1(_03455_),
    .A2(_04024_),
    .ZN(_04408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10083_ (.A1(_02385_),
    .A2(_02396_),
    .ZN(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10084_ (.A1(_04368_),
    .A2(_04409_),
    .ZN(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10085_ (.A1(_02399_),
    .A2(_04168_),
    .ZN(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10086_ (.A1(_04253_),
    .A2(_04410_),
    .B(_04411_),
    .ZN(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10087_ (.A1(\as2650.stack[10][9] ),
    .A2(_04044_),
    .B1(_04046_),
    .B2(\as2650.stack[11][9] ),
    .ZN(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10088_ (.A1(\as2650.stack[9][9] ),
    .A2(_04048_),
    .B1(_04049_),
    .B2(\as2650.stack[8][9] ),
    .ZN(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10089_ (.A1(_04330_),
    .A2(_04413_),
    .A3(_04414_),
    .ZN(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10090_ (.A1(\as2650.stack[13][9] ),
    .A2(_04048_),
    .B1(_04049_),
    .B2(\as2650.stack[12][9] ),
    .ZN(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10091_ (.A1(\as2650.stack[14][9] ),
    .A2(_04044_),
    .B1(_04046_),
    .B2(\as2650.stack[15][9] ),
    .ZN(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10092_ (.A1(_04052_),
    .A2(_04416_),
    .A3(_04417_),
    .ZN(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10093_ (.A1(_04415_),
    .A2(_04418_),
    .Z(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10094_ (.A1(\as2650.stack[5][9] ),
    .A2(_04340_),
    .B1(_04341_),
    .B2(\as2650.stack[4][9] ),
    .ZN(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10095_ (.I(_04420_),
    .ZN(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10096_ (.A1(\as2650.stack[6][9] ),
    .A2(_04338_),
    .B1(_04339_),
    .B2(\as2650.stack[7][9] ),
    .C(_04421_),
    .ZN(_04422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10097_ (.A1(_04375_),
    .A2(_04422_),
    .B(_04061_),
    .ZN(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10098_ (.A1(\as2650.stack[2][9] ),
    .A2(_04116_),
    .B1(_04118_),
    .B2(\as2650.stack[3][9] ),
    .ZN(_04424_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10099_ (.A1(\as2650.stack[1][9] ),
    .A2(_04129_),
    .B1(_04130_),
    .B2(\as2650.stack[0][9] ),
    .ZN(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10100_ (.A1(_04125_),
    .A2(_04424_),
    .A3(_04425_),
    .ZN(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _10101_ (.A1(_03824_),
    .A2(_04419_),
    .B1(_04423_),
    .B2(_04426_),
    .ZN(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10102_ (.A1(_02398_),
    .A2(_04040_),
    .ZN(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10103_ (.A1(_04134_),
    .A2(_04427_),
    .B(_04428_),
    .C(_04236_),
    .ZN(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10104_ (.A1(_04233_),
    .A2(_04412_),
    .B(_04429_),
    .ZN(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10105_ (.A1(_02386_),
    .A2(_04368_),
    .B(_04138_),
    .ZN(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10106_ (.A1(_04013_),
    .A2(_04431_),
    .B(_02396_),
    .ZN(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10107_ (.A1(_04289_),
    .A2(_04430_),
    .B(_04432_),
    .ZN(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10108_ (.I0(_02399_),
    .I1(_04433_),
    .S(_03964_),
    .Z(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10109_ (.A1(_03552_),
    .A2(_04408_),
    .B1(_04434_),
    .B2(_04196_),
    .C(_01680_),
    .ZN(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10110_ (.A1(_04099_),
    .A2(_04433_),
    .B(_03969_),
    .ZN(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10111_ (.A1(_04093_),
    .A2(_04407_),
    .B1(_04435_),
    .B2(_04436_),
    .ZN(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10112_ (.A1(_04406_),
    .A2(_04437_),
    .B(_03717_),
    .ZN(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10113_ (.A1(_01144_),
    .A2(_03875_),
    .B(_04438_),
    .C(_04031_),
    .ZN(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10114_ (.I(_04017_),
    .Z(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10115_ (.A1(\as2650.stack[10][10] ),
    .A2(_04115_),
    .B1(_04117_),
    .B2(\as2650.stack[11][10] ),
    .ZN(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10116_ (.A1(\as2650.stack[9][10] ),
    .A2(_04340_),
    .B1(_04341_),
    .B2(\as2650.stack[8][10] ),
    .ZN(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10117_ (.A1(_03829_),
    .A2(_04440_),
    .A3(_04441_),
    .ZN(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10118_ (.A1(\as2650.stack[13][10] ),
    .A2(_04119_),
    .B1(_04120_),
    .B2(\as2650.stack[12][10] ),
    .ZN(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10119_ (.A1(\as2650.stack[14][10] ),
    .A2(_03989_),
    .B1(_03990_),
    .B2(\as2650.stack[15][10] ),
    .ZN(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10120_ (.A1(_03988_),
    .A2(_04443_),
    .A3(_04444_),
    .ZN(_04445_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10121_ (.A1(_04442_),
    .A2(_04445_),
    .Z(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10122_ (.A1(\as2650.stack[5][10] ),
    .A2(_02478_),
    .B1(_02595_),
    .B2(\as2650.stack[4][10] ),
    .ZN(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10123_ (.I(_04447_),
    .ZN(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10124_ (.A1(\as2650.stack[6][10] ),
    .A2(_04044_),
    .B1(_04046_),
    .B2(\as2650.stack[7][10] ),
    .C(_04448_),
    .ZN(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10125_ (.A1(_04109_),
    .A2(_04449_),
    .B(_03977_),
    .ZN(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10126_ (.I(_02251_),
    .Z(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10127_ (.I(_03834_),
    .Z(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10128_ (.A1(\as2650.stack[2][10] ),
    .A2(_04451_),
    .B1(_04452_),
    .B2(\as2650.stack[3][10] ),
    .ZN(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10129_ (.I(_03979_),
    .Z(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10130_ (.I(_03980_),
    .Z(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10131_ (.A1(\as2650.stack[1][10] ),
    .A2(_04454_),
    .B1(_04455_),
    .B2(\as2650.stack[0][10] ),
    .ZN(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10132_ (.A1(_04330_),
    .A2(_04453_),
    .A3(_04456_),
    .ZN(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _10133_ (.A1(_04257_),
    .A2(_04446_),
    .B1(_04450_),
    .B2(_04457_),
    .ZN(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10134_ (.A1(_03976_),
    .A2(_04458_),
    .ZN(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10135_ (.A1(_03573_),
    .A2(_04173_),
    .B(_04459_),
    .C(_04236_),
    .ZN(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10136_ (.A1(_02410_),
    .A2(_04410_),
    .Z(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10137_ (.A1(_03699_),
    .A2(_04461_),
    .B(_03971_),
    .ZN(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10138_ (.A1(_03573_),
    .A2(_04138_),
    .B(_04462_),
    .ZN(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10139_ (.A1(_04460_),
    .A2(_04463_),
    .ZN(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10140_ (.A1(_03970_),
    .A2(_04464_),
    .ZN(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10141_ (.A1(_02410_),
    .A2(_04165_),
    .B(_04465_),
    .ZN(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10142_ (.A1(_03964_),
    .A2(_02413_),
    .Z(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10143_ (.A1(_04149_),
    .A2(_04466_),
    .B(_04467_),
    .ZN(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10144_ (.A1(_03564_),
    .A2(_03880_),
    .B1(_04468_),
    .B2(_04148_),
    .ZN(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10145_ (.A1(_04439_),
    .A2(_04469_),
    .ZN(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10146_ (.A1(_04154_),
    .A2(_04466_),
    .B(_04398_),
    .ZN(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10147_ (.A1(_04151_),
    .A2(_02413_),
    .ZN(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10148_ (.A1(_04096_),
    .A2(_04472_),
    .Z(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10149_ (.A1(_04470_),
    .A2(_04471_),
    .B1(_04473_),
    .B2(_03650_),
    .ZN(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10150_ (.I(_03809_),
    .Z(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10151_ (.A1(_03428_),
    .A2(_04404_),
    .B(_03814_),
    .ZN(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10152_ (.A1(_04475_),
    .A2(_04476_),
    .B(_03817_),
    .ZN(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10153_ (.A1(\as2650.instruction_args_latch[10] ),
    .A2(_04158_),
    .B1(_04474_),
    .B2(_04477_),
    .ZN(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10154_ (.A1(_03775_),
    .A2(_04478_),
    .ZN(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10155_ (.A1(\as2650.stack[2][11] ),
    .A2(_04451_),
    .B1(_04452_),
    .B2(\as2650.stack[3][11] ),
    .ZN(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10156_ (.A1(\as2650.stack[1][11] ),
    .A2(_04454_),
    .B1(_04455_),
    .B2(\as2650.stack[0][11] ),
    .ZN(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10157_ (.A1(_03830_),
    .A2(_04479_),
    .A3(_04480_),
    .ZN(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10158_ (.A1(\as2650.stack[5][11] ),
    .A2(_04454_),
    .B1(_04455_),
    .B2(\as2650.stack[4][11] ),
    .ZN(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10159_ (.A1(\as2650.stack[6][11] ),
    .A2(_04451_),
    .B1(_04452_),
    .B2(\as2650.stack[7][11] ),
    .ZN(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10160_ (.A1(_04109_),
    .A2(_04482_),
    .A3(_04483_),
    .ZN(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10161_ (.A1(_04481_),
    .A2(_04484_),
    .ZN(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10162_ (.A1(\as2650.stack[10][11] ),
    .A2(_04451_),
    .B1(_04452_),
    .B2(\as2650.stack[11][11] ),
    .ZN(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10163_ (.A1(\as2650.stack[9][11] ),
    .A2(_04454_),
    .B1(_04455_),
    .B2(\as2650.stack[8][11] ),
    .ZN(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10164_ (.A1(_04330_),
    .A2(_04486_),
    .A3(_04487_),
    .ZN(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10165_ (.A1(\as2650.stack[13][11] ),
    .A2(_02479_),
    .B1(_02596_),
    .B2(\as2650.stack[12][11] ),
    .ZN(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10166_ (.A1(\as2650.stack[14][11] ),
    .A2(_02252_),
    .B1(_03835_),
    .B2(\as2650.stack[15][11] ),
    .ZN(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10167_ (.A1(_04109_),
    .A2(_04489_),
    .A3(_04490_),
    .ZN(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10168_ (.A1(_04488_),
    .A2(_04491_),
    .ZN(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10169_ (.I0(_04485_),
    .I1(_04492_),
    .S(_04257_),
    .Z(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10170_ (.A1(_04173_),
    .A2(_04493_),
    .ZN(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10171_ (.A1(_02422_),
    .A2(_03820_),
    .B(_04494_),
    .ZN(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10172_ (.A1(\as2650.PC[10] ),
    .A2(_04410_),
    .ZN(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10173_ (.A1(_02423_),
    .A2(_04496_),
    .B(_02830_),
    .ZN(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10174_ (.A1(_02422_),
    .A2(_04169_),
    .B(_04233_),
    .ZN(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10175_ (.A1(_03641_),
    .A2(_04495_),
    .B1(_04497_),
    .B2(_04498_),
    .ZN(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10176_ (.A1(_03700_),
    .A2(_04496_),
    .B(_03936_),
    .ZN(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _10177_ (.A1(_03622_),
    .A2(_04499_),
    .B1(_04500_),
    .B2(_02419_),
    .ZN(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10178_ (.A1(_03965_),
    .A2(_02422_),
    .ZN(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10179_ (.A1(_04151_),
    .A2(_04501_),
    .B(_04502_),
    .ZN(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10180_ (.A1(_03577_),
    .A2(_04408_),
    .B1(_04503_),
    .B2(_04196_),
    .ZN(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10181_ (.A1(_04154_),
    .A2(_04504_),
    .ZN(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10182_ (.A1(_04439_),
    .A2(_04501_),
    .B(_04146_),
    .ZN(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10183_ (.A1(_04097_),
    .A2(_04502_),
    .B(_03650_),
    .ZN(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10184_ (.A1(_04505_),
    .A2(_04506_),
    .B(_04507_),
    .ZN(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10185_ (.A1(_03571_),
    .A2(_04475_),
    .B(_03876_),
    .ZN(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10186_ (.A1(_03571_),
    .A2(_04475_),
    .B(_04509_),
    .ZN(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10187_ (.A1(_03963_),
    .A2(_04510_),
    .ZN(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10188_ (.A1(_03443_),
    .A2(_04161_),
    .B1(_04508_),
    .B2(_04511_),
    .C(_01446_),
    .ZN(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10189_ (.A1(_02440_),
    .A2(_03820_),
    .ZN(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10190_ (.A1(\as2650.stack[2][12] ),
    .A2(_04219_),
    .B1(_04220_),
    .B2(\as2650.stack[3][12] ),
    .ZN(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10191_ (.I(_04340_),
    .Z(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10192_ (.I(_04341_),
    .Z(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10193_ (.A1(\as2650.stack[1][12] ),
    .A2(_04514_),
    .B1(_04515_),
    .B2(\as2650.stack[0][12] ),
    .ZN(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10194_ (.A1(_04212_),
    .A2(_04513_),
    .A3(_04516_),
    .ZN(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10195_ (.A1(\as2650.stack[5][12] ),
    .A2(_04514_),
    .B1(_04515_),
    .B2(\as2650.stack[4][12] ),
    .ZN(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10196_ (.A1(\as2650.stack[6][12] ),
    .A2(_04219_),
    .B1(_04220_),
    .B2(\as2650.stack[7][12] ),
    .ZN(_04519_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10197_ (.A1(_04375_),
    .A2(_04518_),
    .A3(_04519_),
    .ZN(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10198_ (.A1(_04517_),
    .A2(_04520_),
    .ZN(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10199_ (.A1(\as2650.stack[10][12] ),
    .A2(_04338_),
    .B1(_04339_),
    .B2(\as2650.stack[11][12] ),
    .ZN(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10200_ (.A1(\as2650.stack[9][12] ),
    .A2(_04514_),
    .B1(_04515_),
    .B2(\as2650.stack[8][12] ),
    .ZN(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10201_ (.A1(_04212_),
    .A2(_04522_),
    .A3(_04523_),
    .ZN(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10202_ (.A1(\as2650.stack[13][12] ),
    .A2(_04514_),
    .B1(_04515_),
    .B2(\as2650.stack[12][12] ),
    .ZN(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10203_ (.A1(\as2650.stack[14][12] ),
    .A2(_04338_),
    .B1(_04339_),
    .B2(\as2650.stack[15][12] ),
    .ZN(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10204_ (.A1(_04375_),
    .A2(_04525_),
    .A3(_04526_),
    .ZN(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10205_ (.A1(_03824_),
    .A2(_04524_),
    .A3(_04527_),
    .ZN(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _10206_ (.A1(_04101_),
    .A2(_04521_),
    .B(_04528_),
    .ZN(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10207_ (.A1(_04329_),
    .A2(_04529_),
    .B(_03972_),
    .ZN(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10208_ (.A1(_02439_),
    .A2(_03973_),
    .B(_04497_),
    .ZN(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10209_ (.A1(_02437_),
    .A2(_04531_),
    .Z(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10210_ (.A1(_04512_),
    .A2(_04530_),
    .B1(_04532_),
    .B2(_04166_),
    .ZN(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10211_ (.I0(_02437_),
    .I1(_04533_),
    .S(_03970_),
    .Z(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10212_ (.I0(_02441_),
    .I1(_04534_),
    .S(_04151_),
    .Z(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10213_ (.A1(_03584_),
    .A2(_04408_),
    .B1(_04535_),
    .B2(_04163_),
    .C(_04154_),
    .ZN(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10214_ (.A1(_04439_),
    .A2(_04534_),
    .ZN(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10215_ (.A1(_04536_),
    .A2(_04537_),
    .B(_04200_),
    .ZN(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10216_ (.A1(_03571_),
    .A2(_04475_),
    .B(_03490_),
    .ZN(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10217_ (.A1(_03810_),
    .A2(_04539_),
    .B(_03877_),
    .ZN(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _10218_ (.A1(_02441_),
    .A2(_04097_),
    .A3(_04146_),
    .Z(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10219_ (.A1(_04538_),
    .A2(_04540_),
    .A3(_04541_),
    .ZN(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10220_ (.A1(\as2650.instruction_args_latch[12] ),
    .A2(_03747_),
    .B(_04401_),
    .ZN(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10221_ (.A1(_04088_),
    .A2(_04542_),
    .B(_04543_),
    .ZN(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10222_ (.I(_02869_),
    .Z(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10223_ (.I(_04544_),
    .Z(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10224_ (.I(_04545_),
    .Z(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10225_ (.I(_01398_),
    .Z(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10226_ (.A1(_04547_),
    .A2(_02958_),
    .ZN(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10227_ (.I(_04548_),
    .Z(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10228_ (.A1(_03636_),
    .A2(_03938_),
    .ZN(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10229_ (.A1(_01512_),
    .A2(_04550_),
    .Z(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _10230_ (.A1(_03633_),
    .A2(_01393_),
    .A3(_04547_),
    .A4(_02200_),
    .ZN(_04552_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10231_ (.A1(_02865_),
    .A2(_04552_),
    .Z(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10232_ (.I(_04553_),
    .Z(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10233_ (.A1(_04547_),
    .A2(_02868_),
    .ZN(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10234_ (.A1(_04551_),
    .A2(_04554_),
    .A3(_04555_),
    .ZN(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10235_ (.I(_04556_),
    .ZN(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10236_ (.A1(_03621_),
    .A2(_02848_),
    .ZN(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10237_ (.A1(_02228_),
    .A2(_04552_),
    .ZN(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10238_ (.A1(_01399_),
    .A2(_01404_),
    .B(_01382_),
    .ZN(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10239_ (.A1(_03634_),
    .A2(_03702_),
    .A3(_04560_),
    .Z(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _10240_ (.A1(_00791_),
    .A2(_02230_),
    .Z(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _10241_ (.I(_02838_),
    .Z(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _10242_ (.A1(_04563_),
    .A2(_00768_),
    .A3(_01510_),
    .ZN(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10243_ (.A1(_02865_),
    .A2(_04562_),
    .B(_04564_),
    .C(_02231_),
    .ZN(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10244_ (.A1(_04558_),
    .A2(_04559_),
    .A3(_04561_),
    .A4(_04565_),
    .ZN(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10245_ (.I(_04566_),
    .Z(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10246_ (.A1(_03242_),
    .A2(_04549_),
    .B(_04557_),
    .C(_04567_),
    .ZN(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10247_ (.A1(_00791_),
    .A2(_02230_),
    .ZN(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10248_ (.A1(_02865_),
    .A2(_04569_),
    .ZN(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10249_ (.I(_04570_),
    .Z(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10250_ (.A1(_02228_),
    .A2(_04562_),
    .ZN(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10251_ (.A1(_04556_),
    .A2(_04572_),
    .ZN(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10252_ (.A1(_01376_),
    .A2(_04544_),
    .ZN(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10253_ (.I(_04574_),
    .Z(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10254_ (.A1(_03297_),
    .A2(_03305_),
    .ZN(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10255_ (.A1(_03296_),
    .A2(_04576_),
    .ZN(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10256_ (.I(_03294_),
    .ZN(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10257_ (.A1(_04578_),
    .A2(_03295_),
    .ZN(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10258_ (.A1(_03302_),
    .A2(_04579_),
    .B(_03255_),
    .ZN(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10259_ (.I(_04580_),
    .ZN(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10260_ (.A1(_02226_),
    .A2(_04563_),
    .B1(_02840_),
    .B2(_04577_),
    .C(_04581_),
    .ZN(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10261_ (.I(_02931_),
    .Z(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10262_ (.I(_03008_),
    .Z(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10263_ (.A1(_03269_),
    .A2(_04584_),
    .B(_01803_),
    .ZN(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10264_ (.A1(_01803_),
    .A2(_02187_),
    .ZN(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10265_ (.A1(_02895_),
    .A2(_04585_),
    .B1(_04586_),
    .B2(_04584_),
    .ZN(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10266_ (.A1(_02226_),
    .A2(_04583_),
    .B(_04587_),
    .ZN(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10267_ (.A1(_00788_),
    .A2(_01381_),
    .A3(_02997_),
    .ZN(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10268_ (.A1(_02827_),
    .A2(_04589_),
    .ZN(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10269_ (.I(_04590_),
    .Z(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10270_ (.I(_04591_),
    .Z(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10271_ (.A1(net171),
    .A2(_04591_),
    .ZN(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10272_ (.A1(_01458_),
    .A2(_04592_),
    .B(_04593_),
    .ZN(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10273_ (.A1(_04584_),
    .A2(_02895_),
    .A3(_04594_),
    .B(_04575_),
    .ZN(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10274_ (.A1(_04575_),
    .A2(_04582_),
    .B1(_04588_),
    .B2(_04595_),
    .ZN(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10275_ (.A1(_04573_),
    .A2(_04596_),
    .ZN(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10276_ (.A1(_04010_),
    .A2(_04571_),
    .B(_04597_),
    .ZN(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10277_ (.A1(_02227_),
    .A2(_04568_),
    .B1(_04598_),
    .B2(_04567_),
    .ZN(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10278_ (.A1(_03633_),
    .A2(_00707_),
    .A3(_02842_),
    .Z(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10279_ (.I(_04600_),
    .Z(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10280_ (.I(_04601_),
    .Z(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10281_ (.I(_03937_),
    .Z(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10282_ (.I(_04603_),
    .Z(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10283_ (.I(_04604_),
    .Z(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10284_ (.A1(_04605_),
    .A2(_04601_),
    .ZN(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10285_ (.I(_03742_),
    .Z(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10286_ (.A1(_04546_),
    .A2(_04602_),
    .B(_04606_),
    .C(_04607_),
    .ZN(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10287_ (.I(_03739_),
    .Z(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10288_ (.I(_04609_),
    .Z(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10289_ (.I(_03751_),
    .Z(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10290_ (.A1(_02227_),
    .A2(_04611_),
    .ZN(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10291_ (.A1(_04610_),
    .A2(_04611_),
    .B(_04612_),
    .ZN(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10292_ (.I(_02827_),
    .Z(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10293_ (.A1(_04614_),
    .A2(_04601_),
    .ZN(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10294_ (.A1(_04546_),
    .A2(_04582_),
    .ZN(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10295_ (.A1(_04613_),
    .A2(_04615_),
    .B(_04616_),
    .ZN(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10296_ (.A1(_04599_),
    .A2(_04608_),
    .B1(_04617_),
    .B2(_04607_),
    .ZN(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10297_ (.A1(_04546_),
    .A2(_03678_),
    .B(_04618_),
    .ZN(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10298_ (.A1(_02961_),
    .A2(_04616_),
    .B(_04159_),
    .ZN(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10299_ (.A1(_04619_),
    .A2(_04620_),
    .ZN(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _10300_ (.A1(_03633_),
    .A2(_00707_),
    .A3(_02842_),
    .ZN(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10301_ (.I(_04621_),
    .Z(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _10302_ (.I(_04614_),
    .Z(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10303_ (.I(_03742_),
    .Z(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10304_ (.A1(_04623_),
    .A2(_04624_),
    .ZN(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10305_ (.A1(_04622_),
    .A2(_04625_),
    .ZN(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10306_ (.I(_04626_),
    .Z(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10307_ (.A1(_02269_),
    .A2(_03757_),
    .ZN(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10308_ (.A1(_03658_),
    .A2(_02824_),
    .ZN(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10309_ (.A1(_04628_),
    .A2(_04629_),
    .Z(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10310_ (.I(_04572_),
    .Z(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10311_ (.I(_04631_),
    .Z(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10312_ (.I(_04592_),
    .Z(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10313_ (.A1(_04073_),
    .A2(_04632_),
    .B1(_04633_),
    .B2(net182),
    .ZN(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10314_ (.I(_04631_),
    .Z(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10315_ (.A1(_04635_),
    .A2(_04633_),
    .ZN(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10316_ (.A1(_03644_),
    .A2(_04636_),
    .ZN(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10317_ (.A1(_03645_),
    .A2(_04634_),
    .B1(_04637_),
    .B2(_01775_),
    .ZN(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10318_ (.A1(_04627_),
    .A2(_04638_),
    .B(_04401_),
    .ZN(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10319_ (.A1(_04627_),
    .A2(_04630_),
    .B(_04639_),
    .ZN(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10320_ (.A1(_04563_),
    .A2(_02959_),
    .ZN(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10321_ (.A1(_04602_),
    .A2(_04640_),
    .B(_04606_),
    .C(_04624_),
    .ZN(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10322_ (.I(_04567_),
    .ZN(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10323_ (.I(_04642_),
    .Z(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10324_ (.I0(_03297_),
    .I1(_03296_),
    .S(_03311_),
    .Z(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10325_ (.A1(_04563_),
    .A2(_04574_),
    .ZN(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10326_ (.A1(net193),
    .A2(_04592_),
    .ZN(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10327_ (.A1(_01785_),
    .A2(_04592_),
    .B(_04646_),
    .C(_04549_),
    .ZN(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10328_ (.A1(_04644_),
    .A2(_04645_),
    .B(_04647_),
    .ZN(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10329_ (.A1(_04133_),
    .A2(_04635_),
    .B1(_04573_),
    .B2(_04648_),
    .ZN(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10330_ (.A1(_03411_),
    .A2(_04575_),
    .B(_04556_),
    .C(_04642_),
    .ZN(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10331_ (.A1(_04643_),
    .A2(_04649_),
    .B1(_04650_),
    .B2(_02289_),
    .ZN(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10332_ (.I(_04609_),
    .Z(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10333_ (.A1(_03760_),
    .A2(_04652_),
    .ZN(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10334_ (.A1(_02289_),
    .A2(_03760_),
    .B(_04653_),
    .ZN(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10335_ (.A1(_04641_),
    .A2(_04651_),
    .B1(_04654_),
    .B2(_04626_),
    .ZN(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10336_ (.A1(_03678_),
    .A2(_04640_),
    .B(_04655_),
    .ZN(_04656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10337_ (.A1(_04607_),
    .A2(_04622_),
    .ZN(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10338_ (.A1(_03411_),
    .A2(_04545_),
    .ZN(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10339_ (.A1(_02961_),
    .A2(_04657_),
    .B(_04644_),
    .C(_04658_),
    .ZN(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10340_ (.A1(_03620_),
    .A2(_04656_),
    .A3(_04659_),
    .ZN(_00465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10341_ (.A1(_03453_),
    .A2(_04652_),
    .ZN(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10342_ (.A1(_01804_),
    .A2(_03762_),
    .B(_04660_),
    .ZN(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10343_ (.A1(_04188_),
    .A2(_04632_),
    .B1(_04633_),
    .B2(net197),
    .ZN(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10344_ (.A1(_04583_),
    .A2(_04637_),
    .B1(_04662_),
    .B2(_03645_),
    .ZN(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10345_ (.A1(_04627_),
    .A2(_04663_),
    .B(_04401_),
    .ZN(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10346_ (.A1(_04627_),
    .A2(_04661_),
    .B(_04664_),
    .ZN(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10347_ (.I(_01497_),
    .Z(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10348_ (.A1(_04231_),
    .A2(_04571_),
    .ZN(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10349_ (.A1(net198),
    .A2(_04633_),
    .B(_04666_),
    .ZN(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10350_ (.I(_04289_),
    .Z(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10351_ (.I(_04668_),
    .Z(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10352_ (.A1(_04665_),
    .A2(_04637_),
    .B1(_04667_),
    .B2(_04669_),
    .ZN(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10353_ (.A1(_04626_),
    .A2(_04670_),
    .ZN(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10354_ (.A1(_03765_),
    .A2(_04610_),
    .B(_04602_),
    .ZN(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10355_ (.A1(_01479_),
    .A2(_03765_),
    .B(_04625_),
    .C(_04672_),
    .ZN(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10356_ (.A1(_03620_),
    .A2(_04671_),
    .A3(_04673_),
    .ZN(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10357_ (.A1(_03255_),
    .A2(_03175_),
    .B(_03167_),
    .ZN(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _10358_ (.A1(_03158_),
    .A2(_04674_),
    .ZN(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10359_ (.A1(_04658_),
    .A2(_04675_),
    .ZN(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10360_ (.A1(_01412_),
    .A2(_03677_),
    .Z(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10361_ (.I(_03412_),
    .Z(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10362_ (.A1(_01827_),
    .A2(_03668_),
    .B(_04678_),
    .ZN(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10363_ (.A1(_02822_),
    .A2(_04600_),
    .ZN(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10364_ (.A1(_01466_),
    .A2(_04650_),
    .ZN(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10365_ (.A1(\as2650.debug_psl[5] ),
    .A2(_02931_),
    .ZN(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10366_ (.A1(_04583_),
    .A2(_01602_),
    .B(_02895_),
    .C(_04682_),
    .ZN(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10367_ (.A1(_02331_),
    .A2(_04591_),
    .B(_03126_),
    .ZN(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10368_ (.A1(_01826_),
    .A2(_04591_),
    .B(_04684_),
    .ZN(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10369_ (.A1(_03008_),
    .A2(_04685_),
    .ZN(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10370_ (.A1(_04583_),
    .A2(_01630_),
    .B(_04682_),
    .ZN(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10371_ (.A1(_04683_),
    .A2(_04686_),
    .B1(_04687_),
    .B2(_04584_),
    .ZN(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10372_ (.A1(_04645_),
    .A2(_04675_),
    .B1(_04688_),
    .B2(_04575_),
    .ZN(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10373_ (.A1(_04272_),
    .A2(_04631_),
    .B1(_04573_),
    .B2(_04689_),
    .ZN(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10374_ (.A1(_04643_),
    .A2(_04690_),
    .ZN(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10375_ (.A1(_04681_),
    .A2(_04691_),
    .ZN(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10376_ (.I(_04692_),
    .ZN(_04693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10377_ (.A1(_04658_),
    .A2(_04693_),
    .B(_04676_),
    .ZN(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10378_ (.A1(_04601_),
    .A2(_04679_),
    .B1(_04680_),
    .B2(_04694_),
    .ZN(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10379_ (.A1(_02822_),
    .A2(_04621_),
    .ZN(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10380_ (.A1(_01827_),
    .A2(_03768_),
    .A3(_04623_),
    .A4(_04696_),
    .Z(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10381_ (.A1(_04695_),
    .A2(_04697_),
    .B(_04607_),
    .ZN(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10382_ (.A1(_04624_),
    .A2(_04622_),
    .A3(_04694_),
    .ZN(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10383_ (.A1(_04625_),
    .A2(_04693_),
    .A3(_04699_),
    .ZN(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10384_ (.A1(_03678_),
    .A2(_04640_),
    .B1(_04698_),
    .B2(_04700_),
    .ZN(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10385_ (.A1(_04676_),
    .A2(_04677_),
    .B(_04701_),
    .ZN(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10386_ (.A1(_03756_),
    .A2(_04702_),
    .ZN(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10387_ (.A1(_03030_),
    .A2(_03290_),
    .ZN(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10388_ (.A1(_03144_),
    .A2(_03193_),
    .A3(_03238_),
    .ZN(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10389_ (.A1(_02885_),
    .A2(_02888_),
    .A3(_02971_),
    .A4(_02972_),
    .Z(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10390_ (.A1(_03040_),
    .A2(_03091_),
    .A3(_04704_),
    .A4(_04705_),
    .ZN(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _10391_ (.A1(_03672_),
    .A2(_03668_),
    .A3(_03094_),
    .A4(_03433_),
    .ZN(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10392_ (.A1(_03182_),
    .A2(_02977_),
    .A3(_04611_),
    .A4(_04707_),
    .ZN(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10393_ (.A1(_03773_),
    .A2(_04708_),
    .ZN(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10394_ (.A1(_03242_),
    .A2(_03246_),
    .ZN(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10395_ (.A1(_03258_),
    .A2(_03262_),
    .A3(_03265_),
    .B(_04710_),
    .ZN(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _10396_ (.A1(_02946_),
    .A2(_03006_),
    .A3(_03068_),
    .A4(_03116_),
    .Z(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10397_ (.A1(_03175_),
    .A2(_03215_),
    .A3(_04712_),
    .ZN(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10398_ (.A1(_04711_),
    .A2(_04713_),
    .B(_03310_),
    .ZN(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10399_ (.A1(_01459_),
    .A2(_02826_),
    .ZN(_04715_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10400_ (.A1(_02821_),
    .A2(_01375_),
    .A3(_01380_),
    .A4(_02839_),
    .ZN(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10401_ (.A1(_00624_),
    .A2(_03937_),
    .ZN(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10402_ (.A1(_02821_),
    .A2(_01380_),
    .A3(_01511_),
    .ZN(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10403_ (.A1(\as2650.debug_psu[5] ),
    .A2(\as2650.debug_psu[4] ),
    .A3(net253),
    .ZN(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10404_ (.A1(_02529_),
    .A2(_02533_),
    .A3(_04719_),
    .Z(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _10405_ (.A1(_01473_),
    .A2(\as2650.debug_psl[6] ),
    .A3(\as2650.debug_psl[0] ),
    .A4(\as2650.debug_psl[5] ),
    .ZN(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10406_ (.A1(_01775_),
    .A2(_01785_),
    .A3(_02931_),
    .A4(_04721_),
    .Z(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10407_ (.A1(\as2650.debug_psl[7] ),
    .A2(_00912_),
    .Z(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10408_ (.A1(\as2650.debug_psu[7] ),
    .A2(_02826_),
    .A3(_04720_),
    .B1(_04722_),
    .B2(_04723_),
    .ZN(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10409_ (.A1(_04718_),
    .A2(_04724_),
    .B(_04716_),
    .ZN(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _10410_ (.I(_01459_),
    .ZN(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10411_ (.A1(_04726_),
    .A2(_04718_),
    .Z(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10412_ (.A1(_04715_),
    .A2(_04716_),
    .A3(_04717_),
    .B1(_04725_),
    .B2(_04727_),
    .ZN(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10413_ (.A1(_01633_),
    .A2(_01073_),
    .A3(_00919_),
    .ZN(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10414_ (.A1(_01047_),
    .A2(_02900_),
    .A3(_04729_),
    .ZN(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10415_ (.A1(_03217_),
    .A2(_03125_),
    .ZN(_04731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10416_ (.A1(_03126_),
    .A2(_04728_),
    .B1(_04730_),
    .B2(_04731_),
    .ZN(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10417_ (.A1(_02844_),
    .A2(_03312_),
    .ZN(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10418_ (.A1(_02162_),
    .A2(_01556_),
    .A3(_01574_),
    .A4(_04729_),
    .Z(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10419_ (.A1(_02845_),
    .A2(_04732_),
    .B1(_04733_),
    .B2(_04734_),
    .ZN(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10420_ (.A1(_01331_),
    .A2(_01338_),
    .A3(_01342_),
    .ZN(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _10421_ (.A1(net200),
    .A2(_00631_),
    .A3(_00639_),
    .A4(_01325_),
    .ZN(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10422_ (.A1(_04736_),
    .A2(_04737_),
    .B(_00619_),
    .C(_02835_),
    .ZN(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10423_ (.A1(_02912_),
    .A2(_04735_),
    .B(_04738_),
    .ZN(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10424_ (.A1(_04548_),
    .A2(_04739_),
    .ZN(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10425_ (.A1(_04548_),
    .A2(_04714_),
    .B(_04740_),
    .C(_04555_),
    .ZN(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10426_ (.A1(_00631_),
    .A2(_01086_),
    .B1(_01601_),
    .B2(_00639_),
    .ZN(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10427_ (.A1(_02331_),
    .A2(_01616_),
    .ZN(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10428_ (.A1(_00639_),
    .A2(_01601_),
    .B(_04742_),
    .C(_04743_),
    .ZN(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10429_ (.A1(_01073_),
    .A2(_01592_),
    .B(_04744_),
    .ZN(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10430_ (.A1(_02360_),
    .A2(_02898_),
    .ZN(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10431_ (.A1(_00624_),
    .A2(_00981_),
    .B(_04746_),
    .ZN(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10432_ (.A1(_01556_),
    .A2(_01330_),
    .ZN(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10433_ (.A1(_02346_),
    .A2(_03217_),
    .B1(_02187_),
    .B2(_02239_),
    .C(_04748_),
    .ZN(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10434_ (.A1(_01574_),
    .A2(_01338_),
    .B1(_01342_),
    .B2(_01589_),
    .ZN(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10435_ (.A1(_02185_),
    .A2(_01325_),
    .B1(_01331_),
    .B2(_01556_),
    .C(_04750_),
    .ZN(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10436_ (.A1(_00618_),
    .A2(_02162_),
    .ZN(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10437_ (.A1(_01578_),
    .A2(_02291_),
    .ZN(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10438_ (.A1(_04752_),
    .A2(_04753_),
    .ZN(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _10439_ (.A1(_04747_),
    .A2(_04749_),
    .A3(_04751_),
    .A4(_04754_),
    .ZN(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10440_ (.I(_04742_),
    .ZN(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10441_ (.A1(_02185_),
    .A2(_01324_),
    .B1(_01330_),
    .B2(_01048_),
    .ZN(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10442_ (.A1(_04748_),
    .A2(_04757_),
    .ZN(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10443_ (.A1(_04753_),
    .A2(_04758_),
    .ZN(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10444_ (.A1(_04750_),
    .A2(_04759_),
    .ZN(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _10445_ (.A1(_00624_),
    .A2(_00981_),
    .B1(_04756_),
    .B2(_04743_),
    .C1(_04745_),
    .C2(_04760_),
    .ZN(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10446_ (.A1(\as2650.debug_psl[1] ),
    .A2(_04746_),
    .B1(_04747_),
    .B2(_04761_),
    .C(_04752_),
    .ZN(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10447_ (.A1(_02268_),
    .A2(_04752_),
    .B(_04762_),
    .ZN(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10448_ (.A1(_04745_),
    .A2(_04755_),
    .B(_04763_),
    .ZN(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10449_ (.A1(_04547_),
    .A2(_02868_),
    .A3(_04764_),
    .ZN(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _10450_ (.A1(_04553_),
    .A2(_04741_),
    .A3(_04765_),
    .Z(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10451_ (.A1(_02459_),
    .A2(_00622_),
    .ZN(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10452_ (.A1(_00586_),
    .A2(_00622_),
    .ZN(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10453_ (.A1(net176),
    .A2(_00618_),
    .ZN(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10454_ (.A1(_04768_),
    .A2(_04769_),
    .ZN(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10455_ (.A1(net175),
    .A2(net174),
    .A3(_00617_),
    .A4(_00622_),
    .ZN(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10456_ (.A1(_04770_),
    .A2(_04771_),
    .Z(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10457_ (.A1(_04767_),
    .A2(_04772_),
    .ZN(_04773_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10458_ (.A1(net177),
    .A2(_00618_),
    .A3(_04773_),
    .ZN(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10459_ (.A1(_02469_),
    .A2(_02360_),
    .B(_04772_),
    .ZN(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10460_ (.A1(_04774_),
    .A2(_04775_),
    .ZN(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10461_ (.A1(_04770_),
    .A2(_04771_),
    .ZN(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10462_ (.A1(_04772_),
    .A2(_04777_),
    .ZN(_04778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10463_ (.A1(_00595_),
    .A2(_00621_),
    .ZN(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10464_ (.A1(net175),
    .A2(_00617_),
    .A3(_04779_),
    .ZN(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10465_ (.A1(_02434_),
    .A2(_00614_),
    .B1(_02345_),
    .B2(_02451_),
    .ZN(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10466_ (.A1(net175),
    .A2(_00630_),
    .ZN(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10467_ (.A1(_04779_),
    .A2(_04782_),
    .Z(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10468_ (.A1(net173),
    .A2(_00617_),
    .A3(_04783_),
    .ZN(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10469_ (.A1(_04779_),
    .A2(_04782_),
    .B(_04784_),
    .ZN(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10470_ (.A1(_04771_),
    .A2(_04781_),
    .A3(_04785_),
    .ZN(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10471_ (.A1(_04780_),
    .A2(_04786_),
    .Z(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10472_ (.A1(_00587_),
    .A2(net176),
    .A3(_00623_),
    .A4(_00631_),
    .ZN(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10473_ (.A1(_02469_),
    .A2(_01622_),
    .B(_04767_),
    .ZN(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10474_ (.A1(_04788_),
    .A2(_04789_),
    .ZN(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10475_ (.I(_04790_),
    .ZN(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10476_ (.A1(_04780_),
    .A2(_04786_),
    .ZN(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10477_ (.A1(_04787_),
    .A2(_04791_),
    .B(_04792_),
    .ZN(_04793_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10478_ (.A1(_04778_),
    .A2(_04793_),
    .ZN(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10479_ (.A1(_04778_),
    .A2(_04793_),
    .ZN(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10480_ (.A1(_04788_),
    .A2(_04795_),
    .ZN(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10481_ (.A1(_04794_),
    .A2(_04796_),
    .ZN(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10482_ (.A1(_04776_),
    .A2(_04797_),
    .ZN(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10483_ (.A1(_04776_),
    .A2(_04797_),
    .ZN(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10484_ (.A1(_00605_),
    .A2(_00636_),
    .Z(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10485_ (.A1(_00602_),
    .A2(_01340_),
    .ZN(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10486_ (.A1(_00600_),
    .A2(_01336_),
    .ZN(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10487_ (.A1(_04800_),
    .A2(_04801_),
    .A3(_04802_),
    .ZN(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10488_ (.A1(_00595_),
    .A2(_00597_),
    .A3(_01321_),
    .A4(_01327_),
    .Z(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10489_ (.A1(net174),
    .A2(_01321_),
    .B1(_01327_),
    .B2(_00598_),
    .ZN(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10490_ (.A1(_04804_),
    .A2(_04805_),
    .ZN(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10491_ (.A1(_04803_),
    .A2(_04806_),
    .Z(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10492_ (.A1(net173),
    .A2(_01322_),
    .ZN(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10493_ (.A1(_00606_),
    .A2(_01341_),
    .Z(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10494_ (.A1(_00603_),
    .A2(_01335_),
    .ZN(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10495_ (.A1(_00601_),
    .A2(_01327_),
    .ZN(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10496_ (.A1(_04809_),
    .A2(_04810_),
    .A3(_04811_),
    .ZN(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10497_ (.A1(_04808_),
    .A2(_04812_),
    .Z(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10498_ (.A1(_04807_),
    .A2(_04813_),
    .ZN(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10499_ (.A1(_04810_),
    .A2(_04811_),
    .ZN(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10500_ (.A1(_04810_),
    .A2(_04811_),
    .ZN(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10501_ (.A1(_04809_),
    .A2(_04815_),
    .B(_04816_),
    .ZN(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10502_ (.A1(_04807_),
    .A2(_04813_),
    .ZN(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10503_ (.A1(_04817_),
    .A2(_04818_),
    .ZN(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10504_ (.A1(_04804_),
    .A2(_04803_),
    .A3(_04805_),
    .ZN(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10505_ (.A1(_00605_),
    .A2(_00629_),
    .Z(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10506_ (.A1(_00602_),
    .A2(_00636_),
    .ZN(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10507_ (.A1(_00600_),
    .A2(_01340_),
    .ZN(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10508_ (.A1(_04821_),
    .A2(_04822_),
    .A3(_04823_),
    .Z(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10509_ (.I(_04804_),
    .ZN(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10510_ (.I(_00594_),
    .Z(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10511_ (.A1(_04826_),
    .A2(_01326_),
    .ZN(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10512_ (.A1(_00591_),
    .A2(_01321_),
    .ZN(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10513_ (.A1(_00596_),
    .A2(_01335_),
    .ZN(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10514_ (.A1(_04827_),
    .A2(_04828_),
    .A3(_04829_),
    .Z(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10515_ (.A1(_04825_),
    .A2(_04830_),
    .Z(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10516_ (.A1(_04824_),
    .A2(_04831_),
    .Z(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10517_ (.A1(_04801_),
    .A2(_04802_),
    .ZN(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10518_ (.A1(_04801_),
    .A2(_04802_),
    .ZN(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10519_ (.A1(_04800_),
    .A2(_04833_),
    .B(_04834_),
    .ZN(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10520_ (.A1(_04820_),
    .A2(_04832_),
    .A3(_04835_),
    .ZN(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10521_ (.A1(_04814_),
    .A2(_04819_),
    .B(_04836_),
    .ZN(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10522_ (.A1(_04825_),
    .A2(_04830_),
    .ZN(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10523_ (.A1(_04824_),
    .A2(_04831_),
    .B(_04838_),
    .ZN(_04839_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10524_ (.A1(_04827_),
    .A2(_04828_),
    .Z(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10525_ (.A1(_04827_),
    .A2(_04828_),
    .Z(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10526_ (.A1(_04829_),
    .A2(_04840_),
    .B(_04841_),
    .ZN(_04842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10527_ (.A1(_00595_),
    .A2(_01335_),
    .ZN(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10528_ (.A1(_00592_),
    .A2(_01326_),
    .ZN(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10529_ (.A1(_00598_),
    .A2(_01340_),
    .ZN(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10530_ (.A1(_04843_),
    .A2(_04844_),
    .A3(_04845_),
    .ZN(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10531_ (.A1(_00606_),
    .A2(_00620_),
    .ZN(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10532_ (.A1(_00603_),
    .A2(_00630_),
    .ZN(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10533_ (.A1(_00601_),
    .A2(_00637_),
    .ZN(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10534_ (.A1(_04847_),
    .A2(_04848_),
    .A3(_04849_),
    .Z(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10535_ (.A1(_04842_),
    .A2(_04846_),
    .A3(_04850_),
    .Z(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10536_ (.A1(_04822_),
    .A2(_04823_),
    .ZN(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10537_ (.A1(_04822_),
    .A2(_04823_),
    .ZN(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10538_ (.A1(_04821_),
    .A2(_04852_),
    .B(_04853_),
    .ZN(_04854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10539_ (.A1(_00588_),
    .A2(_01322_),
    .ZN(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10540_ (.A1(_04854_),
    .A2(_04855_),
    .Z(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10541_ (.A1(_04854_),
    .A2(_04855_),
    .ZN(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10542_ (.A1(_04856_),
    .A2(_04857_),
    .ZN(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10543_ (.A1(_04839_),
    .A2(_04851_),
    .A3(_04858_),
    .ZN(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10544_ (.A1(_04820_),
    .A2(_04832_),
    .ZN(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10545_ (.A1(_04820_),
    .A2(_04832_),
    .ZN(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10546_ (.A1(_04835_),
    .A2(_04860_),
    .B(_04861_),
    .ZN(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10547_ (.A1(_04859_),
    .A2(_04862_),
    .ZN(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10548_ (.A1(_04817_),
    .A2(_04818_),
    .Z(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10549_ (.A1(_00607_),
    .A2(_01337_),
    .ZN(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10550_ (.A1(_00604_),
    .A2(_01328_),
    .ZN(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10551_ (.A1(net172),
    .A2(_01323_),
    .ZN(_04867_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10552_ (.A1(_04866_),
    .A2(_04867_),
    .Z(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10553_ (.A1(_04866_),
    .A2(_04867_),
    .Z(_04869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10554_ (.A1(_04865_),
    .A2(_04868_),
    .B(_04869_),
    .ZN(_04870_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10555_ (.A1(_04808_),
    .A2(_04812_),
    .Z(_04871_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10556_ (.A1(_04870_),
    .A2(_04871_),
    .Z(_04872_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10557_ (.A1(_04866_),
    .A2(_04867_),
    .A3(_04865_),
    .Z(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10558_ (.A1(net203),
    .A2(_00607_),
    .A3(_01323_),
    .A4(_01329_),
    .ZN(_04874_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10559_ (.A1(_04873_),
    .A2(_04874_),
    .ZN(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10560_ (.A1(_04872_),
    .A2(_04875_),
    .Z(_04876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10561_ (.A1(_04864_),
    .A2(_04876_),
    .ZN(_04877_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _10562_ (.A1(_04836_),
    .A2(_04814_),
    .A3(_04819_),
    .Z(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10563_ (.A1(_04837_),
    .A2(_04878_),
    .Z(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10564_ (.A1(_04870_),
    .A2(_04871_),
    .Z(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10565_ (.A1(_04864_),
    .A2(_04880_),
    .ZN(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10566_ (.A1(_04879_),
    .A2(_04881_),
    .Z(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10567_ (.A1(_04879_),
    .A2(_04864_),
    .A3(_04880_),
    .ZN(_04883_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10568_ (.A1(_04877_),
    .A2(_04882_),
    .B(_04883_),
    .ZN(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10569_ (.A1(_04837_),
    .A2(_04863_),
    .Z(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10570_ (.A1(_04884_),
    .A2(_04885_),
    .ZN(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10571_ (.A1(_04837_),
    .A2(_04863_),
    .B(_04886_),
    .ZN(_04887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10572_ (.A1(_04859_),
    .A2(_04862_),
    .ZN(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10573_ (.A1(_04839_),
    .A2(_04851_),
    .Z(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10574_ (.A1(_04839_),
    .A2(_04851_),
    .Z(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10575_ (.A1(_04858_),
    .A2(_04889_),
    .B(_04890_),
    .ZN(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10576_ (.A1(_04842_),
    .A2(_04846_),
    .ZN(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10577_ (.A1(_04842_),
    .A2(_04846_),
    .ZN(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10578_ (.A1(_04850_),
    .A2(_04892_),
    .B(_04893_),
    .ZN(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10579_ (.A1(_00606_),
    .A2(_00616_),
    .ZN(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10580_ (.A1(_00603_),
    .A2(_00620_),
    .ZN(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10581_ (.A1(_00599_),
    .A2(_00629_),
    .ZN(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10582_ (.A1(_04896_),
    .A2(_04897_),
    .ZN(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10583_ (.A1(_04895_),
    .A2(_04898_),
    .ZN(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10584_ (.A1(_04843_),
    .A2(_04844_),
    .Z(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10585_ (.A1(_04843_),
    .A2(_04844_),
    .Z(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10586_ (.A1(_04845_),
    .A2(_04900_),
    .B(_04901_),
    .ZN(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10587_ (.A1(_04826_),
    .A2(_01339_),
    .ZN(_04903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10588_ (.A1(_00592_),
    .A2(_01334_),
    .ZN(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10589_ (.A1(_00597_),
    .A2(_00637_),
    .ZN(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10590_ (.A1(_04903_),
    .A2(_04904_),
    .A3(_04905_),
    .ZN(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10591_ (.A1(_04902_),
    .A2(_04906_),
    .ZN(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10592_ (.A1(_04899_),
    .A2(_04907_),
    .Z(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10593_ (.A1(_00588_),
    .A2(_01328_),
    .ZN(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10594_ (.A1(_04848_),
    .A2(_04849_),
    .Z(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10595_ (.A1(_04848_),
    .A2(_04849_),
    .Z(_04911_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10596_ (.A1(_04847_),
    .A2(_04910_),
    .B(_04911_),
    .ZN(_04912_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10597_ (.A1(_00584_),
    .A2(_01322_),
    .ZN(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10598_ (.A1(_04912_),
    .A2(_04913_),
    .ZN(_04914_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10599_ (.A1(_04909_),
    .A2(_04914_),
    .Z(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10600_ (.A1(_04894_),
    .A2(_04908_),
    .A3(_04915_),
    .ZN(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10601_ (.A1(_04856_),
    .A2(_04891_),
    .A3(_04916_),
    .Z(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10602_ (.A1(_04888_),
    .A2(_04917_),
    .ZN(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10603_ (.I(_04918_),
    .ZN(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10604_ (.A1(_04888_),
    .A2(_04917_),
    .ZN(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10605_ (.A1(_04887_),
    .A2(_04919_),
    .B(_04920_),
    .ZN(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10606_ (.A1(_04891_),
    .A2(_04916_),
    .ZN(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10607_ (.A1(_04891_),
    .A2(_04916_),
    .ZN(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10608_ (.A1(_04856_),
    .A2(_04922_),
    .B(_04923_),
    .ZN(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10609_ (.A1(_00586_),
    .A2(_01324_),
    .A3(_04912_),
    .ZN(_04925_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10610_ (.A1(_02459_),
    .A2(_01329_),
    .A3(_04914_),
    .ZN(_04926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10611_ (.A1(_04925_),
    .A2(_04926_),
    .ZN(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10612_ (.A1(_04894_),
    .A2(_04908_),
    .ZN(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10613_ (.A1(_04894_),
    .A2(_04908_),
    .ZN(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10614_ (.A1(_04915_),
    .A2(_04928_),
    .B(_04929_),
    .ZN(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10615_ (.A1(_04902_),
    .A2(_04906_),
    .ZN(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10616_ (.A1(_04899_),
    .A2(_04907_),
    .B(_04931_),
    .ZN(_04932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10617_ (.A1(_00600_),
    .A2(_00621_),
    .ZN(_04933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10618_ (.A1(_00604_),
    .A2(_00615_),
    .ZN(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10619_ (.A1(_04933_),
    .A2(_04934_),
    .ZN(_04935_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10620_ (.A1(_04903_),
    .A2(_04904_),
    .Z(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10621_ (.A1(_04903_),
    .A2(_04904_),
    .Z(_04937_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10622_ (.A1(_04905_),
    .A2(_04936_),
    .B(_04937_),
    .ZN(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10623_ (.A1(_02450_),
    .A2(_02433_),
    .A3(_00634_),
    .A4(_01591_),
    .ZN(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10624_ (.A1(_04826_),
    .A2(_00635_),
    .B1(_01339_),
    .B2(_00591_),
    .ZN(_04940_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10625_ (.A1(_04939_),
    .A2(_04940_),
    .ZN(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10626_ (.A1(_00596_),
    .A2(_00629_),
    .ZN(_04942_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10627_ (.I(_04942_),
    .ZN(_04943_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10628_ (.A1(_04941_),
    .A2(_04943_),
    .Z(_04944_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10629_ (.A1(_04938_),
    .A2(_04944_),
    .ZN(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10630_ (.A1(_04935_),
    .A2(_04945_),
    .Z(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10631_ (.A1(_04932_),
    .A2(_04946_),
    .Z(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10632_ (.A1(_00589_),
    .A2(_01336_),
    .ZN(_04948_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _10633_ (.A1(_02393_),
    .A2(_02345_),
    .A3(_04897_),
    .B1(_04898_),
    .B2(_04895_),
    .ZN(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10634_ (.A1(_00584_),
    .A2(_01328_),
    .ZN(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10635_ (.A1(_04949_),
    .A2(_04950_),
    .ZN(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10636_ (.A1(_04948_),
    .A2(_04951_),
    .ZN(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10637_ (.A1(_04947_),
    .A2(_04952_),
    .Z(_04953_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10638_ (.A1(_04930_),
    .A2(_04953_),
    .Z(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10639_ (.A1(_04927_),
    .A2(_04954_),
    .Z(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10640_ (.A1(_04924_),
    .A2(_04955_),
    .ZN(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10641_ (.A1(_04924_),
    .A2(_04955_),
    .ZN(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10642_ (.A1(_04921_),
    .A2(_04956_),
    .B(_04957_),
    .ZN(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10643_ (.A1(_04930_),
    .A2(_04953_),
    .Z(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10644_ (.A1(_04927_),
    .A2(_04954_),
    .B(_04959_),
    .ZN(_04960_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10645_ (.A1(_00587_),
    .A2(_01330_),
    .A3(_04949_),
    .ZN(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10646_ (.A1(net176),
    .A2(_01337_),
    .A3(_04951_),
    .ZN(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10647_ (.A1(_04961_),
    .A2(_04962_),
    .ZN(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10648_ (.A1(_04932_),
    .A2(_04946_),
    .ZN(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10649_ (.A1(_04947_),
    .A2(_04952_),
    .ZN(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10650_ (.A1(_04964_),
    .A2(_04965_),
    .ZN(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10651_ (.A1(_04938_),
    .A2(_04944_),
    .ZN(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10652_ (.A1(_04935_),
    .A2(_04945_),
    .B(_04967_),
    .ZN(_04968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10653_ (.A1(_00601_),
    .A2(_00616_),
    .ZN(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10654_ (.A1(_04941_),
    .A2(_04943_),
    .B(_04939_),
    .ZN(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10655_ (.A1(_02450_),
    .A2(_02434_),
    .A3(_00627_),
    .A4(_00634_),
    .ZN(_04971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10656_ (.A1(_04826_),
    .A2(_00628_),
    .B1(_00636_),
    .B2(_00592_),
    .ZN(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10657_ (.A1(_04971_),
    .A2(_04972_),
    .Z(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10658_ (.A1(_00597_),
    .A2(_00620_),
    .ZN(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10659_ (.A1(_04973_),
    .A2(_04974_),
    .ZN(_04975_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10660_ (.A1(_04970_),
    .A2(_04975_),
    .ZN(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10661_ (.A1(_04969_),
    .A2(_04976_),
    .Z(_04977_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10662_ (.A1(_04968_),
    .A2(_04977_),
    .Z(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10663_ (.A1(_04933_),
    .A2(_04934_),
    .ZN(_04979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10664_ (.A1(_00588_),
    .A2(_01341_),
    .ZN(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10665_ (.A1(_00585_),
    .A2(_01336_),
    .ZN(_04981_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10666_ (.A1(_04979_),
    .A2(_04980_),
    .A3(_04981_),
    .Z(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10667_ (.A1(_04978_),
    .A2(_04982_),
    .Z(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10668_ (.A1(_04966_),
    .A2(_04983_),
    .Z(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10669_ (.A1(_04963_),
    .A2(_04984_),
    .ZN(_04985_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10670_ (.A1(_04960_),
    .A2(_04985_),
    .Z(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10671_ (.A1(_04960_),
    .A2(_04985_),
    .ZN(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10672_ (.A1(_04958_),
    .A2(_04986_),
    .B(_04987_),
    .ZN(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10673_ (.A1(_04966_),
    .A2(_04983_),
    .Z(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10674_ (.A1(_04963_),
    .A2(_04984_),
    .B(_04989_),
    .ZN(_04990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10675_ (.A1(net177),
    .A2(_01337_),
    .B(_04979_),
    .ZN(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10676_ (.A1(_00587_),
    .A2(_01338_),
    .A3(_04979_),
    .ZN(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10677_ (.A1(_04980_),
    .A2(_04991_),
    .B(_04992_),
    .ZN(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10678_ (.A1(_04968_),
    .A2(_04977_),
    .ZN(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10679_ (.A1(_04978_),
    .A2(_04982_),
    .ZN(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10680_ (.A1(_04994_),
    .A2(_04995_),
    .ZN(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10681_ (.A1(_04973_),
    .A2(_04974_),
    .ZN(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10682_ (.A1(_04971_),
    .A2(_04997_),
    .ZN(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10683_ (.A1(_00598_),
    .A2(_00616_),
    .ZN(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10684_ (.A1(_04783_),
    .A2(_04999_),
    .Z(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10685_ (.A1(_04998_),
    .A2(_05000_),
    .Z(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _10686_ (.A1(_02406_),
    .A2(_01644_),
    .A3(_04976_),
    .B1(_04975_),
    .B2(_04970_),
    .ZN(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10687_ (.A1(_05001_),
    .A2(_05002_),
    .Z(_05003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10688_ (.A1(_00589_),
    .A2(_00637_),
    .ZN(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10689_ (.A1(_00585_),
    .A2(_01341_),
    .ZN(_05005_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10690_ (.A1(_05004_),
    .A2(_05005_),
    .Z(_05006_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10691_ (.A1(_05003_),
    .A2(_05006_),
    .Z(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10692_ (.A1(_04996_),
    .A2(_05007_),
    .Z(_05008_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10693_ (.A1(_04993_),
    .A2(_05008_),
    .ZN(_05009_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10694_ (.A1(_04990_),
    .A2(_05009_),
    .Z(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10695_ (.A1(_04990_),
    .A2(_05009_),
    .ZN(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10696_ (.A1(_05010_),
    .A2(_05011_),
    .ZN(_05012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10697_ (.A1(_04988_),
    .A2(_05012_),
    .B(_05010_),
    .ZN(_05013_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10698_ (.A1(_04996_),
    .A2(_05007_),
    .Z(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10699_ (.A1(_04993_),
    .A2(_05008_),
    .B(_05014_),
    .ZN(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10700_ (.A1(_05004_),
    .A2(_05005_),
    .Z(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10701_ (.A1(_05001_),
    .A2(_05002_),
    .ZN(_05017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10702_ (.A1(_05003_),
    .A2(_05006_),
    .ZN(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10703_ (.A1(_05017_),
    .A2(_05018_),
    .ZN(_05019_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10704_ (.A1(_00586_),
    .A2(_02459_),
    .A3(_00630_),
    .A4(_00638_),
    .ZN(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10705_ (.A1(_02460_),
    .A2(_00627_),
    .B1(_02317_),
    .B2(_02468_),
    .ZN(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10706_ (.A1(_05020_),
    .A2(_05021_),
    .ZN(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10707_ (.A1(_04998_),
    .A2(_05000_),
    .Z(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10708_ (.A1(_04771_),
    .A2(_04781_),
    .ZN(_05024_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10709_ (.A1(_05024_),
    .A2(_04785_),
    .Z(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10710_ (.A1(_05023_),
    .A2(_05025_),
    .ZN(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10711_ (.A1(_05022_),
    .A2(_05026_),
    .Z(_05027_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10712_ (.A1(_05019_),
    .A2(_05027_),
    .Z(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10713_ (.A1(_05016_),
    .A2(_05028_),
    .Z(_05029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10714_ (.A1(_05015_),
    .A2(_05029_),
    .ZN(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10715_ (.A1(_05015_),
    .A2(_05029_),
    .ZN(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10716_ (.A1(_05013_),
    .A2(_05030_),
    .B(_05031_),
    .ZN(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10717_ (.I(_05028_),
    .ZN(_05033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10718_ (.A1(_05019_),
    .A2(_05027_),
    .ZN(_05034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10719_ (.A1(_05016_),
    .A2(_05033_),
    .B(_05034_),
    .ZN(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _10720_ (.A1(_04998_),
    .A2(_05000_),
    .A3(_05025_),
    .B1(_05022_),
    .B2(_05026_),
    .ZN(_05036_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10721_ (.A1(_04787_),
    .A2(_04791_),
    .Z(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10722_ (.A1(_05036_),
    .A2(_05037_),
    .ZN(_05038_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10723_ (.A1(_05020_),
    .A2(_05038_),
    .Z(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10724_ (.A1(_05035_),
    .A2(_05039_),
    .ZN(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10725_ (.A1(_05035_),
    .A2(_05039_),
    .ZN(_05041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10726_ (.A1(_05032_),
    .A2(_05040_),
    .B(_05041_),
    .ZN(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10727_ (.A1(_05020_),
    .A2(_05038_),
    .ZN(_05043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10728_ (.A1(_05036_),
    .A2(_05037_),
    .B(_05043_),
    .ZN(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10729_ (.A1(_04788_),
    .A2(_04795_),
    .Z(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10730_ (.I(_05045_),
    .ZN(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10731_ (.A1(_05044_),
    .A2(_05046_),
    .ZN(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10732_ (.A1(_05044_),
    .A2(_05046_),
    .ZN(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10733_ (.A1(_05042_),
    .A2(_05047_),
    .B(_05048_),
    .ZN(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10734_ (.A1(_04799_),
    .A2(_05049_),
    .ZN(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10735_ (.A1(_04553_),
    .A2(_04774_),
    .ZN(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _10736_ (.A1(_04798_),
    .A2(_05050_),
    .A3(_05051_),
    .ZN(_05052_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10737_ (.A1(_04799_),
    .A2(_05049_),
    .ZN(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10738_ (.A1(_05044_),
    .A2(_05045_),
    .A3(_05042_),
    .Z(_05054_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10739_ (.A1(_05035_),
    .A2(_05039_),
    .A3(_05032_),
    .Z(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _10740_ (.A1(_05015_),
    .A2(_05029_),
    .A3(_05013_),
    .Z(_05056_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10741_ (.A1(_04988_),
    .A2(_05012_),
    .Z(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10742_ (.A1(_04958_),
    .A2(_04986_),
    .Z(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _10743_ (.A1(_04921_),
    .A2(_04956_),
    .ZN(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10744_ (.A1(_04887_),
    .A2(_04918_),
    .Z(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _10745_ (.A1(_04884_),
    .A2(_04885_),
    .ZN(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10746_ (.A1(_04877_),
    .A2(_04882_),
    .Z(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10747_ (.A1(_04880_),
    .A2(_04876_),
    .ZN(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _10748_ (.A1(_04864_),
    .A2(_05063_),
    .ZN(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10749_ (.A1(_04872_),
    .A2(_04875_),
    .Z(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10750_ (.A1(_04873_),
    .A2(_04874_),
    .Z(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10751_ (.A1(net203),
    .A2(_01324_),
    .B1(_01331_),
    .B2(net202),
    .ZN(_05067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10752_ (.A1(_02376_),
    .A2(_02239_),
    .B(_05067_),
    .ZN(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10753_ (.A1(_05066_),
    .A2(_05068_),
    .Z(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10754_ (.A1(_05062_),
    .A2(_05064_),
    .A3(_05065_),
    .A4(_05069_),
    .ZN(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10755_ (.A1(_05059_),
    .A2(_05060_),
    .A3(_05061_),
    .A4(_05070_),
    .ZN(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10756_ (.A1(_05056_),
    .A2(_05057_),
    .A3(_05058_),
    .A4(_05071_),
    .ZN(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10757_ (.A1(_05053_),
    .A2(_05054_),
    .A3(_05055_),
    .A4(_05072_),
    .ZN(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10758_ (.A1(_04551_),
    .A2(_04570_),
    .Z(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10759_ (.A1(_05052_),
    .A2(_05073_),
    .B(_05074_),
    .ZN(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10760_ (.A1(_04304_),
    .A2(_04572_),
    .ZN(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10761_ (.A1(_04766_),
    .A2(_05075_),
    .B(_05076_),
    .ZN(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10762_ (.A1(_04566_),
    .A2(_04550_),
    .B(_04726_),
    .ZN(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10763_ (.A1(_04567_),
    .A2(_05077_),
    .B(_05078_),
    .ZN(_05079_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _10764_ (.A1(_01412_),
    .A2(_03679_),
    .A3(_02864_),
    .Z(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10765_ (.I(_05080_),
    .ZN(_05081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10766_ (.I(_02868_),
    .Z(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10767_ (.A1(_01412_),
    .A2(_02960_),
    .ZN(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10768_ (.A1(_05082_),
    .A2(_02959_),
    .B(_05083_),
    .ZN(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10769_ (.A1(_05079_),
    .A2(_05081_),
    .B(_05084_),
    .ZN(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10770_ (.A1(_01803_),
    .A2(_02829_),
    .ZN(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10771_ (.A1(_01880_),
    .A2(_04605_),
    .B(_03452_),
    .ZN(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10772_ (.I(_02827_),
    .Z(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10773_ (.A1(_02269_),
    .A2(_05088_),
    .ZN(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10774_ (.A1(_01859_),
    .A2(_04603_),
    .B(_02976_),
    .ZN(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10775_ (.A1(net164),
    .A2(_04604_),
    .ZN(_05091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10776_ (.A1(_01460_),
    .A2(_02828_),
    .B(_03240_),
    .ZN(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10777_ (.A1(_05089_),
    .A2(_05090_),
    .B1(_05091_),
    .B2(_05092_),
    .ZN(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10778_ (.A1(_01896_),
    .A2(_04604_),
    .ZN(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10779_ (.A1(_01826_),
    .A2(_02828_),
    .B(_03196_),
    .ZN(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10780_ (.A1(_02226_),
    .A2(_05088_),
    .ZN(_05096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10781_ (.A1(_01847_),
    .A2(_00820_),
    .B(_03751_),
    .ZN(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10782_ (.A1(_05094_),
    .A2(_05095_),
    .B1(_05096_),
    .B2(_05097_),
    .ZN(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10783_ (.A1(\as2650.debug_psu[7] ),
    .A2(_02826_),
    .B(_04723_),
    .ZN(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10784_ (.A1(\as2650.debug_psl[2] ),
    .A2(_05088_),
    .ZN(_05100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10785_ (.A1(_01866_),
    .A2(_04603_),
    .B(_03042_),
    .ZN(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10786_ (.A1(_03675_),
    .A2(_05099_),
    .B1(_05100_),
    .B2(_05101_),
    .ZN(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10787_ (.A1(_05093_),
    .A2(_05098_),
    .A3(_05102_),
    .ZN(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10788_ (.A1(_01475_),
    .A2(_04614_),
    .ZN(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10789_ (.A1(_03470_),
    .A2(_05104_),
    .ZN(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10790_ (.A1(\as2650.debug_psu[4] ),
    .A2(_04605_),
    .B(_05105_),
    .ZN(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10791_ (.A1(_05086_),
    .A2(_05087_),
    .B(_05103_),
    .C(_05106_),
    .ZN(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10792_ (.A1(_05088_),
    .A2(_05079_),
    .ZN(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10793_ (.A1(_04726_),
    .A2(_03671_),
    .A3(_04604_),
    .ZN(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10794_ (.A1(_05108_),
    .A2(_05109_),
    .B(_04696_),
    .ZN(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10795_ (.A1(_02163_),
    .A2(_03738_),
    .ZN(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_2 _10796_ (.A1(_03093_),
    .A2(_01590_),
    .B1(_01576_),
    .B2(_03433_),
    .C1(_02891_),
    .C2(_02904_),
    .ZN(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10797_ (.A1(_03658_),
    .A2(_01557_),
    .B1(_01602_),
    .B2(_03469_),
    .ZN(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10798_ (.A1(_01669_),
    .A2(_03269_),
    .B1(_03218_),
    .B2(_03240_),
    .C(_05113_),
    .ZN(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10799_ (.A1(_03668_),
    .A2(_03146_),
    .B(_05114_),
    .ZN(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10800_ (.A1(_05111_),
    .A2(_05112_),
    .A3(_05115_),
    .B(_05082_),
    .ZN(_05116_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10801_ (.A1(_04544_),
    .A2(_05079_),
    .A3(_05116_),
    .ZN(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10802_ (.A1(_04544_),
    .A2(_04714_),
    .ZN(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10803_ (.A1(_05111_),
    .A2(_05118_),
    .B(_05116_),
    .ZN(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _10804_ (.A1(_03667_),
    .A2(_01625_),
    .B1(_01638_),
    .B2(_03243_),
    .ZN(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10805_ (.A1(_03469_),
    .A2(_01609_),
    .B1(_01625_),
    .B2(_03667_),
    .C(_05120_),
    .ZN(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10806_ (.A1(_03674_),
    .A2(_01647_),
    .Z(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10807_ (.A1(_03093_),
    .A2(_01596_),
    .B1(_01609_),
    .B2(_03469_),
    .ZN(_05123_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10808_ (.I(_05123_),
    .ZN(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10809_ (.A1(_01581_),
    .A2(_01582_),
    .ZN(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10810_ (.A1(_01575_),
    .A2(_01563_),
    .B(_05125_),
    .ZN(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10811_ (.A1(_03093_),
    .A2(_01596_),
    .ZN(_05127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10812_ (.A1(_01369_),
    .A2(_05126_),
    .B(_05127_),
    .ZN(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10813_ (.A1(_03042_),
    .A2(_05126_),
    .ZN(_05129_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10814_ (.I(_01550_),
    .ZN(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10815_ (.A1(_03750_),
    .A2(_05130_),
    .B1(_01568_),
    .B2(_02975_),
    .ZN(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10816_ (.A1(_02976_),
    .A2(_01568_),
    .ZN(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10817_ (.A1(_02891_),
    .A2(_01550_),
    .B(_05132_),
    .ZN(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10818_ (.A1(_05129_),
    .A2(_05131_),
    .A3(_05133_),
    .ZN(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10819_ (.A1(_03243_),
    .A2(_01638_),
    .B(_05128_),
    .C(_05134_),
    .ZN(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10820_ (.A1(_05121_),
    .A2(_05122_),
    .A3(_05124_),
    .A4(_05135_),
    .Z(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10821_ (.A1(_05082_),
    .A2(_05136_),
    .ZN(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10822_ (.A1(_03674_),
    .A2(_01647_),
    .Z(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10823_ (.A1(_05131_),
    .A2(_05132_),
    .Z(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10824_ (.A1(_05129_),
    .A2(_05139_),
    .B(_05128_),
    .ZN(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10825_ (.A1(_05123_),
    .A2(_05140_),
    .ZN(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10826_ (.A1(_03470_),
    .A2(_01609_),
    .B1(_01625_),
    .B2(_03667_),
    .C(_05141_),
    .ZN(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10827_ (.A1(_03671_),
    .A2(_01638_),
    .ZN(_05143_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10828_ (.A1(_05120_),
    .A2(_05142_),
    .B(_05143_),
    .ZN(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10829_ (.A1(_02268_),
    .A2(_03674_),
    .A3(_01647_),
    .ZN(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10830_ (.A1(_02268_),
    .A2(_05138_),
    .B1(_05122_),
    .B2(_05144_),
    .C(_05145_),
    .ZN(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10831_ (.A1(_05137_),
    .A2(_05146_),
    .ZN(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10832_ (.A1(_04680_),
    .A2(_05147_),
    .ZN(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10833_ (.A1(_01459_),
    .A2(_03671_),
    .B(_02828_),
    .ZN(_05149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10834_ (.A1(_03739_),
    .A2(_05149_),
    .B(_04600_),
    .ZN(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10835_ (.A1(_05117_),
    .A2(_05119_),
    .A3(_05148_),
    .B1(_05150_),
    .B2(_05108_),
    .ZN(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10836_ (.A1(_05110_),
    .A2(_05151_),
    .ZN(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10837_ (.A1(_03740_),
    .A2(_05152_),
    .ZN(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10838_ (.A1(_03740_),
    .A2(_05107_),
    .B(_05153_),
    .C(_05080_),
    .ZN(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10839_ (.A1(_05118_),
    .A2(_05147_),
    .ZN(_05155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10840_ (.A1(_05085_),
    .A2(_05154_),
    .B1(_05155_),
    .B2(_04677_),
    .C(_02978_),
    .ZN(_05156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10841_ (.A1(_02978_),
    .A2(_04709_),
    .B(_05156_),
    .ZN(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10842_ (.A1(_04703_),
    .A2(_04706_),
    .B1(_05157_),
    .B2(_03030_),
    .ZN(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10843_ (.A1(_03756_),
    .A2(_05158_),
    .ZN(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10844_ (.I(_05146_),
    .ZN(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10845_ (.A1(_04545_),
    .A2(_03329_),
    .B1(_05137_),
    .B2(_05159_),
    .ZN(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10846_ (.A1(_03636_),
    .A2(_03938_),
    .A3(_04643_),
    .ZN(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10847_ (.A1(_03311_),
    .A2(_04549_),
    .ZN(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10848_ (.A1(_03937_),
    .A2(_04589_),
    .ZN(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10849_ (.A1(\as2650.debug_psl[7] ),
    .A2(_04718_),
    .ZN(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10850_ (.A1(_04718_),
    .A2(_05099_),
    .B(_05164_),
    .C(_04716_),
    .ZN(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10851_ (.A1(_00619_),
    .A2(_04590_),
    .B1(_05163_),
    .B2(_01467_),
    .C(_05165_),
    .ZN(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10852_ (.A1(_03126_),
    .A2(_05166_),
    .B(_04731_),
    .ZN(_05167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10853_ (.A1(_03008_),
    .A2(_05167_),
    .B(_04733_),
    .ZN(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10854_ (.A1(_02912_),
    .A2(_05168_),
    .ZN(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10855_ (.A1(net201),
    .A2(_02912_),
    .B(_04574_),
    .C(_05169_),
    .ZN(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10856_ (.A1(_05162_),
    .A2(_05170_),
    .B(_04555_),
    .ZN(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10857_ (.A1(_04555_),
    .A2(_04763_),
    .B(_05171_),
    .C(_04554_),
    .ZN(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10858_ (.A1(_05074_),
    .A2(_05052_),
    .A3(_05172_),
    .B1(_04631_),
    .B2(_04349_),
    .ZN(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10859_ (.A1(_01467_),
    .A2(_05161_),
    .B1(_05173_),
    .B2(_04643_),
    .ZN(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10860_ (.A1(_05082_),
    .A2(_02959_),
    .A3(_04615_),
    .A4(_05111_),
    .ZN(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10861_ (.A1(_03291_),
    .A2(_03739_),
    .ZN(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10862_ (.A1(_01467_),
    .A2(_03291_),
    .B(_05176_),
    .ZN(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10863_ (.A1(_04615_),
    .A2(_05177_),
    .B(_05160_),
    .ZN(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10864_ (.A1(_05080_),
    .A2(_05178_),
    .ZN(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10865_ (.A1(_05174_),
    .A2(_05175_),
    .B(_05179_),
    .ZN(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10866_ (.A1(_05080_),
    .A2(_05174_),
    .ZN(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10867_ (.A1(_03740_),
    .A2(_05180_),
    .B(_05181_),
    .ZN(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10868_ (.A1(_05083_),
    .A2(_05160_),
    .B1(_05182_),
    .B2(_05084_),
    .ZN(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10869_ (.A1(_02860_),
    .A2(_05183_),
    .B(_03292_),
    .ZN(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10870_ (.A1(_03371_),
    .A2(_04703_),
    .A3(_05184_),
    .ZN(_00470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10871_ (.A1(_04089_),
    .A2(_03869_),
    .B(_02214_),
    .ZN(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10872_ (.A1(_03963_),
    .A2(_05185_),
    .B(_01849_),
    .ZN(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _10873_ (.A1(_02829_),
    .A2(_04621_),
    .ZN(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10874_ (.A1(_01848_),
    .A2(_04611_),
    .ZN(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10875_ (.A1(_04610_),
    .A2(_03752_),
    .B(_05188_),
    .ZN(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10876_ (.A1(_02214_),
    .A2(_04024_),
    .ZN(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10877_ (.A1(_05187_),
    .A2(_05189_),
    .B(_05190_),
    .ZN(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10878_ (.A1(_04624_),
    .A2(_05187_),
    .ZN(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10879_ (.A1(_04329_),
    .A2(_04569_),
    .ZN(_05193_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10880_ (.A1(_02231_),
    .A2(_05193_),
    .ZN(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10881_ (.I(_05163_),
    .Z(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10882_ (.I(_05195_),
    .Z(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10883_ (.I(_05163_),
    .Z(_05197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10884_ (.A1(_01848_),
    .A2(_05197_),
    .ZN(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10885_ (.A1(_02239_),
    .A2(_05196_),
    .B(_05198_),
    .ZN(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10886_ (.A1(_05194_),
    .A2(_05199_),
    .Z(_05200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10887_ (.A1(_03644_),
    .A2(_05200_),
    .ZN(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10888_ (.A1(_01849_),
    .A2(_03697_),
    .B(_05192_),
    .C(_05201_),
    .ZN(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10889_ (.A1(_02214_),
    .A2(_03818_),
    .ZN(_05203_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10890_ (.A1(_03716_),
    .A2(_05203_),
    .ZN(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10891_ (.A1(_01681_),
    .A2(_05191_),
    .B(_05202_),
    .C(_05204_),
    .ZN(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10892_ (.A1(_01450_),
    .A2(_05186_),
    .A3(_05205_),
    .Z(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10893_ (.I(_05206_),
    .Z(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10894_ (.I(_05204_),
    .Z(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10895_ (.A1(_02254_),
    .A2(_03857_),
    .ZN(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _10896_ (.A1(_04623_),
    .A2(_01663_),
    .A3(_03741_),
    .ZN(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10897_ (.A1(_01860_),
    .A2(_02977_),
    .ZN(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10898_ (.A1(_04602_),
    .A2(_04629_),
    .A3(_05209_),
    .A4(_05210_),
    .ZN(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10899_ (.A1(_02148_),
    .A2(_02216_),
    .A3(_05208_),
    .B(_05211_),
    .ZN(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10900_ (.A1(_04162_),
    .A2(_05212_),
    .ZN(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10901_ (.A1(_05187_),
    .A2(_05190_),
    .B(_04099_),
    .ZN(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10902_ (.I(_03635_),
    .Z(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10903_ (.A1(_01859_),
    .A2(_05197_),
    .ZN(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10904_ (.A1(_01564_),
    .A2(_05197_),
    .B(_05216_),
    .ZN(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10905_ (.A1(_02197_),
    .A2(_05215_),
    .ZN(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10906_ (.A1(_05215_),
    .A2(_05217_),
    .B1(_05218_),
    .B2(_01859_),
    .ZN(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10907_ (.I(_04569_),
    .Z(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10908_ (.A1(_05208_),
    .A2(_05193_),
    .B1(_05219_),
    .B2(_05220_),
    .ZN(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10909_ (.A1(_02483_),
    .A2(_05221_),
    .Z(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10910_ (.A1(_02257_),
    .A2(_05208_),
    .B(_05222_),
    .C(_03697_),
    .ZN(_05223_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10911_ (.A1(_02475_),
    .A2(_03753_),
    .B(_05214_),
    .C(_05223_),
    .ZN(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10912_ (.A1(_05213_),
    .A2(_05224_),
    .ZN(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10913_ (.I(_01433_),
    .Z(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10914_ (.A1(_05208_),
    .A2(_05207_),
    .B(_05226_),
    .ZN(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10915_ (.A1(_05207_),
    .A2(_05225_),
    .B(_05227_),
    .ZN(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10916_ (.A1(_01866_),
    .A2(_03856_),
    .Z(_05228_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10917_ (.A1(_02247_),
    .A2(_03660_),
    .ZN(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10918_ (.A1(_02216_),
    .A2(_05228_),
    .Z(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10919_ (.A1(_04606_),
    .A2(_04653_),
    .A3(_05229_),
    .B1(_05230_),
    .B2(_02148_),
    .ZN(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10920_ (.A1(_02257_),
    .A2(_05228_),
    .ZN(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10921_ (.A1(_01866_),
    .A2(_05195_),
    .ZN(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10922_ (.A1(_02291_),
    .A2(_05195_),
    .B(_05233_),
    .ZN(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10923_ (.A1(_01867_),
    .A2(_05218_),
    .B1(_05234_),
    .B2(_05215_),
    .ZN(_05235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10924_ (.A1(_03862_),
    .A2(_05193_),
    .B1(_05235_),
    .B2(_05220_),
    .ZN(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10925_ (.A1(_02483_),
    .A2(_05236_),
    .ZN(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10926_ (.A1(_05232_),
    .A2(_05237_),
    .B(_04668_),
    .ZN(_05238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10927_ (.A1(_01869_),
    .A2(_03631_),
    .B(_05238_),
    .ZN(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10928_ (.A1(_04439_),
    .A2(_05231_),
    .B1(_05239_),
    .B2(_05214_),
    .C(_05203_),
    .ZN(_05240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10929_ (.A1(_05203_),
    .A2(_05228_),
    .B(_05240_),
    .C(_04161_),
    .ZN(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10930_ (.A1(_03776_),
    .A2(_05230_),
    .B(_04159_),
    .ZN(_05242_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10931_ (.A1(_05241_),
    .A2(_05242_),
    .ZN(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10932_ (.A1(_01881_),
    .A2(_03453_),
    .B(_04622_),
    .C(_04660_),
    .ZN(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10933_ (.A1(_01867_),
    .A2(_02254_),
    .ZN(_05244_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10934_ (.A1(_02530_),
    .A2(_05244_),
    .Z(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10935_ (.A1(_02148_),
    .A2(_02216_),
    .A3(_05245_),
    .ZN(_05246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10936_ (.A1(_05209_),
    .A2(_05243_),
    .B(_05246_),
    .ZN(_05247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10937_ (.A1(_01879_),
    .A2(_05195_),
    .ZN(_05248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10938_ (.A1(_01592_),
    .A2(_05197_),
    .B(_05248_),
    .ZN(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10939_ (.A1(_01879_),
    .A2(_05218_),
    .B1(_05249_),
    .B2(_05215_),
    .ZN(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10940_ (.A1(_04100_),
    .A2(_05220_),
    .B(_03825_),
    .ZN(_05251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10941_ (.A1(_05220_),
    .A2(_05250_),
    .B(_05251_),
    .ZN(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10942_ (.A1(_02483_),
    .A2(_05252_),
    .Z(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10943_ (.A1(_02257_),
    .A2(_05245_),
    .B(_05253_),
    .C(_03631_),
    .ZN(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10944_ (.A1(_02531_),
    .A2(_03645_),
    .B(_05214_),
    .C(_05254_),
    .ZN(_05255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10945_ (.A1(_01681_),
    .A2(_05247_),
    .B(_05255_),
    .ZN(_05256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10946_ (.A1(_05207_),
    .A2(_05245_),
    .B(_05226_),
    .ZN(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10947_ (.A1(_05207_),
    .A2(_05256_),
    .B(_05257_),
    .ZN(_00474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10948_ (.I(_05192_),
    .Z(_05258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10949_ (.I(_05196_),
    .Z(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10950_ (.A1(_04632_),
    .A2(_05259_),
    .B(_03622_),
    .ZN(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10951_ (.A1(_04529_),
    .A2(_04635_),
    .B1(_05259_),
    .B2(net198),
    .ZN(_05261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10952_ (.A1(_04669_),
    .A2(_05261_),
    .ZN(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10953_ (.A1(_01888_),
    .A2(_05260_),
    .B(_05262_),
    .ZN(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _10954_ (.I(_01888_),
    .ZN(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10955_ (.A1(_05264_),
    .A2(_03663_),
    .B(_05209_),
    .ZN(_05265_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10956_ (.A1(_04672_),
    .A2(_05265_),
    .ZN(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10957_ (.A1(_05258_),
    .A2(_05263_),
    .B1(_05266_),
    .B2(_04162_),
    .C(_01446_),
    .ZN(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10958_ (.I(_01896_),
    .ZN(_05267_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10959_ (.A1(_01365_),
    .A2(_04100_),
    .B1(_05196_),
    .B2(net199),
    .ZN(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10960_ (.A1(_05267_),
    .A2(_05196_),
    .B1(_05268_),
    .B2(_04668_),
    .ZN(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10961_ (.A1(_04668_),
    .A2(_03866_),
    .A3(_04571_),
    .ZN(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _10962_ (.A1(_01897_),
    .A2(_03631_),
    .B1(_04571_),
    .B2(_05269_),
    .C(_05270_),
    .ZN(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10963_ (.A1(_03669_),
    .A2(_02824_),
    .ZN(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10964_ (.A1(_05267_),
    .A2(_03669_),
    .B(_05187_),
    .C(_05272_),
    .ZN(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10965_ (.A1(_05258_),
    .A2(_05271_),
    .ZN(_05274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10966_ (.A1(_01440_),
    .A2(_05273_),
    .B(_05274_),
    .ZN(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10967_ (.A1(_03614_),
    .A2(_05271_),
    .B(_05275_),
    .C(_03718_),
    .ZN(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10968_ (.A1(_03896_),
    .A2(_04632_),
    .B1(_05259_),
    .B2(net200),
    .ZN(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10969_ (.A1(_04669_),
    .A2(_05276_),
    .ZN(_05277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10970_ (.A1(_01903_),
    .A2(_05260_),
    .B(_05277_),
    .ZN(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10971_ (.A1(_03771_),
    .A2(_04610_),
    .ZN(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10972_ (.A1(_01903_),
    .A2(_03771_),
    .B(_05192_),
    .C(_05279_),
    .ZN(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10973_ (.A1(_05258_),
    .A2(_05278_),
    .B(_05280_),
    .C(_04031_),
    .ZN(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10974_ (.A1(_03919_),
    .A2(_04635_),
    .B1(_05259_),
    .B2(net201),
    .ZN(_05281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10975_ (.A1(_04669_),
    .A2(_05281_),
    .ZN(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10976_ (.A1(net29),
    .A2(_05260_),
    .B(_05282_),
    .ZN(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10977_ (.A1(_01910_),
    .A2(_03773_),
    .B(_05176_),
    .C(_05192_),
    .ZN(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10978_ (.I(_03619_),
    .Z(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10979_ (.A1(_05258_),
    .A2(_05283_),
    .B(_05284_),
    .C(_05285_),
    .ZN(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10980_ (.A1(_01448_),
    .A2(_03713_),
    .ZN(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10981_ (.I(_05286_),
    .Z(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10982_ (.I0(net36),
    .I1(\as2650.irqs_latch[1] ),
    .S(_05287_),
    .Z(_05288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10983_ (.I(_05288_),
    .Z(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10984_ (.A1(net37),
    .A2(_05287_),
    .ZN(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10985_ (.A1(_01273_),
    .A2(_05287_),
    .B(_05289_),
    .ZN(_00480_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10986_ (.I0(net38),
    .I1(\as2650.irqs_latch[3] ),
    .S(_05287_),
    .Z(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10987_ (.I(_05290_),
    .Z(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10988_ (.I(_05286_),
    .Z(_05291_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10989_ (.I0(\as2650.trap ),
    .I1(\as2650.irqs_latch[4] ),
    .S(_05291_),
    .Z(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10990_ (.I(_05292_),
    .Z(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10991_ (.I0(net39),
    .I1(\as2650.irqs_latch[5] ),
    .S(_05291_),
    .Z(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10992_ (.I(_05293_),
    .Z(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10993_ (.I0(net40),
    .I1(\as2650.irqs_latch[6] ),
    .S(_05291_),
    .Z(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10994_ (.I(_05294_),
    .Z(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10995_ (.I0(net41),
    .I1(\as2650.irqs_latch[7] ),
    .S(_05291_),
    .Z(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10996_ (.I(_05295_),
    .Z(_00485_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10997_ (.I(_04559_),
    .ZN(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10998_ (.A1(_02229_),
    .A2(_04558_),
    .A3(_04564_),
    .ZN(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10999_ (.A1(_04558_),
    .A2(_05296_),
    .B1(_05297_),
    .B2(\as2650.trap ),
    .ZN(_05298_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11000_ (.A1(_03756_),
    .A2(_05298_),
    .ZN(_00486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11001_ (.I(_03728_),
    .Z(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11002_ (.I(_05299_),
    .Z(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11003_ (.I(_03729_),
    .Z(_05301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11004_ (.A1(net131),
    .A2(_05301_),
    .B(_05226_),
    .ZN(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11005_ (.A1(_02904_),
    .A2(_05300_),
    .B(_05302_),
    .ZN(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11006_ (.A1(net132),
    .A2(_05301_),
    .B(_05226_),
    .ZN(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11007_ (.A1(_01558_),
    .A2(_05300_),
    .B(_05303_),
    .ZN(_00488_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11008_ (.I(_03729_),
    .Z(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11009_ (.I(_01433_),
    .Z(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11010_ (.A1(net133),
    .A2(_05304_),
    .B(_05305_),
    .ZN(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11011_ (.A1(_01576_),
    .A2(_05300_),
    .B(_05306_),
    .ZN(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11012_ (.A1(net134),
    .A2(_05304_),
    .B(_05305_),
    .ZN(_05307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11013_ (.A1(_01590_),
    .A2(_05300_),
    .B(_05307_),
    .ZN(_00490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11014_ (.I(_05299_),
    .Z(_05308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11015_ (.A1(net135),
    .A2(_05304_),
    .B(_05305_),
    .ZN(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11016_ (.A1(_01603_),
    .A2(_05308_),
    .B(_05309_),
    .ZN(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11017_ (.A1(net136),
    .A2(_05304_),
    .B(_05305_),
    .ZN(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11018_ (.A1(_03146_),
    .A2(_05308_),
    .B(_05310_),
    .ZN(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11019_ (.A1(net137),
    .A2(_05299_),
    .B(_01434_),
    .ZN(_05311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11020_ (.A1(_01630_),
    .A2(_05308_),
    .B(_05311_),
    .ZN(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11021_ (.A1(net138),
    .A2(_05299_),
    .B(_01434_),
    .ZN(_05312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11022_ (.A1(_02162_),
    .A2(_05308_),
    .B(_05312_),
    .ZN(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11023_ (.A1(_00645_),
    .A2(_03706_),
    .B(net130),
    .ZN(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11024_ (.A1(_03727_),
    .A2(_05301_),
    .A3(_05313_),
    .ZN(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11025_ (.I(_03743_),
    .Z(_05314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11026_ (.I(_05314_),
    .Z(_05315_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11027_ (.A1(net124),
    .A2(_03744_),
    .ZN(_05316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11028_ (.A1(_03752_),
    .A2(_05315_),
    .B(_05316_),
    .C(_05285_),
    .ZN(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11029_ (.A1(net125),
    .A2(_03744_),
    .ZN(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11030_ (.A1(_03757_),
    .A2(_05315_),
    .B(_05317_),
    .C(_05285_),
    .ZN(_00497_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11031_ (.A1(net126),
    .A2(_03744_),
    .ZN(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11032_ (.A1(_03760_),
    .A2(_05315_),
    .B(_05318_),
    .C(_05285_),
    .ZN(_00498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11033_ (.I(_05314_),
    .Z(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11034_ (.A1(net127),
    .A2(_05319_),
    .ZN(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11035_ (.I(_03619_),
    .Z(_05321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11036_ (.A1(_03762_),
    .A2(_05315_),
    .B(_05320_),
    .C(_05321_),
    .ZN(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11037_ (.I(_05314_),
    .Z(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11038_ (.A1(net128),
    .A2(_05319_),
    .ZN(_05323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11039_ (.A1(_03765_),
    .A2(_05322_),
    .B(_05323_),
    .C(_05321_),
    .ZN(_00500_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11040_ (.A1(net129),
    .A2(_05319_),
    .ZN(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11041_ (.A1(_03768_),
    .A2(_05322_),
    .B(_05324_),
    .C(_05321_),
    .ZN(_00501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11042_ (.A1(\as2650.ext_io_addr[6] ),
    .A2(_05319_),
    .ZN(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11043_ (.A1(_03771_),
    .A2(_05322_),
    .B(_05325_),
    .C(_05321_),
    .ZN(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11044_ (.A1(\as2650.ext_io_addr[7] ),
    .A2(_05314_),
    .ZN(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11045_ (.A1(_03773_),
    .A2(_05322_),
    .B(_05326_),
    .C(_03620_),
    .ZN(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11046_ (.A1(\as2650.io_bus_we ),
    .A2(_03729_),
    .ZN(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11047_ (.A1(_01359_),
    .A2(_05301_),
    .B(_05327_),
    .C(_03727_),
    .ZN(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11048_ (.A1(_01517_),
    .A2(_00375_),
    .A3(_01528_),
    .Z(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11049_ (.I(_05328_),
    .Z(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11050_ (.A1(_00669_),
    .A2(_01434_),
    .ZN(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _11051_ (.A1(_03613_),
    .A2(_02201_),
    .A3(_03590_),
    .A4(_04678_),
    .ZN(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _11052_ (.A1(_03369_),
    .A2(_02938_),
    .A3(_03393_),
    .A4(_05330_),
    .ZN(_05331_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11053_ (.A1(_02010_),
    .A2(_03588_),
    .B1(_05329_),
    .B2(_05331_),
    .ZN(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11054_ (.A1(_01477_),
    .A2(_04652_),
    .ZN(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11055_ (.A1(_02150_),
    .A2(_02874_),
    .A3(_02877_),
    .ZN(_05333_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _11056_ (.A1(_05333_),
    .A2(_02852_),
    .A3(_02862_),
    .A4(_02871_),
    .Z(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11057_ (.I(_05334_),
    .Z(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _11058_ (.A1(_04614_),
    .A2(_05335_),
    .ZN(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11059_ (.A1(_05332_),
    .A2(_05336_),
    .ZN(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11060_ (.I(_05337_),
    .Z(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11061_ (.I(_01476_),
    .Z(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11062_ (.A1(_04605_),
    .A2(_02962_),
    .ZN(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _11063_ (.A1(_05339_),
    .A2(_04609_),
    .A3(_05340_),
    .ZN(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11064_ (.I(_05341_),
    .Z(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11065_ (.I(_01353_),
    .Z(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11066_ (.A1(_05332_),
    .A2(_05336_),
    .B(_05341_),
    .C(_05343_),
    .ZN(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11067_ (.I(_05344_),
    .Z(_05345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11068_ (.A1(_02957_),
    .A2(_05342_),
    .B1(_05345_),
    .B2(\as2650.regs[2][0] ),
    .ZN(_05346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11069_ (.A1(_02956_),
    .A2(_05338_),
    .B(_05346_),
    .ZN(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11070_ (.I(_03007_),
    .Z(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11071_ (.A1(_05347_),
    .A2(_05342_),
    .B1(_05345_),
    .B2(\as2650.regs[2][1] ),
    .ZN(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11072_ (.A1(_03035_),
    .A2(_05338_),
    .B(_05348_),
    .ZN(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11073_ (.I(_03069_),
    .Z(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11074_ (.A1(_05349_),
    .A2(_05342_),
    .B1(_05345_),
    .B2(\as2650.regs[2][2] ),
    .ZN(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11075_ (.A1(_03088_),
    .A2(_05338_),
    .B(_05350_),
    .ZN(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11076_ (.I(_03117_),
    .Z(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11077_ (.A1(_05351_),
    .A2(_05342_),
    .B1(_05345_),
    .B2(\as2650.regs[2][3] ),
    .ZN(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11078_ (.A1(_03138_),
    .A2(_05338_),
    .B(_05352_),
    .ZN(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11079_ (.I(_05337_),
    .Z(_05353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11080_ (.I(_03176_),
    .Z(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11081_ (.I(_05341_),
    .Z(_05355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11082_ (.I(_05344_),
    .Z(_05356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11083_ (.A1(_05354_),
    .A2(_05355_),
    .B1(_05356_),
    .B2(\as2650.regs[2][4] ),
    .ZN(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11084_ (.A1(_03188_),
    .A2(_05353_),
    .B(_05357_),
    .ZN(_00511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11085_ (.I(_03216_),
    .Z(_05358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11086_ (.A1(_05358_),
    .A2(_05355_),
    .B1(_05356_),
    .B2(\as2650.regs[2][5] ),
    .ZN(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11087_ (.A1(_03233_),
    .A2(_05353_),
    .B(_05359_),
    .ZN(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11088_ (.I(_03267_),
    .Z(_05360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11089_ (.A1(_05360_),
    .A2(_05355_),
    .B1(_05356_),
    .B2(\as2650.regs[2][6] ),
    .ZN(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11090_ (.A1(_03285_),
    .A2(_05353_),
    .B(_05361_),
    .ZN(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11091_ (.I(_03329_),
    .Z(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11092_ (.A1(_05362_),
    .A2(_05355_),
    .B1(_05356_),
    .B2(\as2650.regs[2][7] ),
    .ZN(_05363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11093_ (.A1(_03328_),
    .A2(_05353_),
    .B(_05363_),
    .ZN(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11094_ (.A1(_01477_),
    .A2(_04652_),
    .A3(_05336_),
    .ZN(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11095_ (.I(_05364_),
    .Z(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11096_ (.A1(_01813_),
    .A2(_01353_),
    .ZN(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11097_ (.I(_05366_),
    .Z(_05367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11098_ (.A1(_01002_),
    .A2(_05367_),
    .ZN(_05368_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11099_ (.A1(_02228_),
    .A2(_02261_),
    .ZN(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11100_ (.I(_05369_),
    .Z(_05370_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11101_ (.A1(_03412_),
    .A2(_02256_),
    .A3(_05370_),
    .ZN(_05371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11102_ (.A1(_04564_),
    .A2(_04562_),
    .B(_05370_),
    .ZN(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11103_ (.I(_05372_),
    .Z(_05373_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _11104_ (.A1(_02822_),
    .A2(_04603_),
    .A3(_02256_),
    .A4(_05370_),
    .ZN(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11105_ (.A1(_02235_),
    .A2(_04560_),
    .A3(_04548_),
    .Z(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11106_ (.I(_05375_),
    .Z(_05376_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11107_ (.A1(_01513_),
    .A2(_02484_),
    .Z(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11108_ (.A1(_02235_),
    .A2(_04554_),
    .Z(_05378_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _11109_ (.A1(_05376_),
    .A2(_05377_),
    .A3(_05378_),
    .ZN(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _11110_ (.A1(_05371_),
    .A2(_05373_),
    .A3(_05374_),
    .A4(_05379_),
    .ZN(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11111_ (.A1(_01477_),
    .A2(_05380_),
    .ZN(_05381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11112_ (.I(_05381_),
    .Z(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11113_ (.A1(_02955_),
    .A2(_05365_),
    .B(_05368_),
    .C(_05382_),
    .ZN(_05383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11114_ (.A1(_01813_),
    .A2(_01431_),
    .ZN(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11115_ (.A1(_01393_),
    .A2(_01634_),
    .ZN(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11116_ (.A1(_04545_),
    .A2(_03677_),
    .A3(_05385_),
    .ZN(_05386_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11117_ (.A1(_05384_),
    .A2(_05386_),
    .Z(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11118_ (.I(_05387_),
    .Z(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11119_ (.A1(_02484_),
    .A2(_04560_),
    .A3(_04549_),
    .ZN(_05389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11120_ (.A1(_01513_),
    .A2(_02234_),
    .ZN(_05390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11121_ (.I(_05390_),
    .Z(_05391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11122_ (.A1(_02235_),
    .A2(_04554_),
    .ZN(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11123_ (.I(_05392_),
    .Z(_05393_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11124_ (.A1(_05391_),
    .A2(_05393_),
    .A3(_05372_),
    .A4(_05374_),
    .Z(_05394_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11125_ (.A1(_05389_),
    .A2(_05371_),
    .A3(_05394_),
    .ZN(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11126_ (.A1(_05339_),
    .A2(_05395_),
    .Z(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11127_ (.I(_05396_),
    .Z(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11128_ (.I(_05374_),
    .Z(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11129_ (.I(_05398_),
    .Z(_05399_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11130_ (.A1(_03412_),
    .A2(_02256_),
    .A3(_05370_),
    .Z(_05400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11131_ (.I(_05400_),
    .Z(_05401_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11132_ (.I(_05376_),
    .Z(_05402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11133_ (.I(_05390_),
    .Z(_05403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11134_ (.I(_05392_),
    .Z(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11135_ (.A1(_04562_),
    .A2(_05369_),
    .ZN(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11136_ (.I(_05405_),
    .Z(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11137_ (.I(_05405_),
    .Z(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11138_ (.A1(net202),
    .A2(_05407_),
    .ZN(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11139_ (.A1(_04010_),
    .A2(_05406_),
    .B(_05408_),
    .C(_05391_),
    .ZN(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11140_ (.A1(\as2650.chirpchar[0] ),
    .A2(_05403_),
    .B(_05404_),
    .C(_05409_),
    .ZN(_05410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11141_ (.I(_05378_),
    .Z(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11142_ (.A1(net202),
    .A2(net171),
    .A3(_05411_),
    .ZN(_05412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11143_ (.I(_05375_),
    .Z(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11144_ (.A1(_05410_),
    .A2(_05412_),
    .B(_05413_),
    .ZN(_05414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11145_ (.A1(_02947_),
    .A2(_05402_),
    .B(_05414_),
    .ZN(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11146_ (.I(_05400_),
    .Z(_05416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11147_ (.A1(_02227_),
    .A2(_05416_),
    .ZN(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11148_ (.I(_05398_),
    .Z(_05418_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11149_ (.A1(_05401_),
    .A2(_05415_),
    .B(_05417_),
    .C(_05418_),
    .ZN(_05419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11150_ (.A1(_01849_),
    .A2(_05399_),
    .B(_05419_),
    .ZN(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11151_ (.A1(_05397_),
    .A2(_05420_),
    .ZN(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11152_ (.A1(_05383_),
    .A2(_05388_),
    .A3(_05421_),
    .ZN(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11153_ (.A1(_05384_),
    .A2(_05386_),
    .ZN(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11154_ (.I(_05423_),
    .Z(_05424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11155_ (.I(_01497_),
    .Z(_05425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11156_ (.I(_02823_),
    .Z(_05426_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _11157_ (.A1(_05425_),
    .A2(_05426_),
    .A3(_04623_),
    .A4(_05335_),
    .ZN(_05427_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _11158_ (.A1(_05427_),
    .A2(_05396_),
    .A3(_05384_),
    .A4(_05423_),
    .ZN(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11159_ (.I(_05428_),
    .Z(_05429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11160_ (.A1(_02957_),
    .A2(_05424_),
    .B1(_05429_),
    .B2(\as2650.regs[4][0] ),
    .ZN(_05430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11161_ (.A1(_05422_),
    .A2(_05430_),
    .ZN(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11162_ (.A1(_02973_),
    .A2(_03033_),
    .Z(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11163_ (.I(_05366_),
    .Z(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11164_ (.A1(_05431_),
    .A2(_05427_),
    .B1(_05432_),
    .B2(_01020_),
    .C(_05396_),
    .ZN(_05433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11165_ (.I(_05371_),
    .Z(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11166_ (.I(_05434_),
    .Z(_05435_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11167_ (.I(_04874_),
    .ZN(_05436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11168_ (.I(_05378_),
    .Z(_05437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11169_ (.A1(_05436_),
    .A2(_05067_),
    .B(_05437_),
    .ZN(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11170_ (.A1(_04073_),
    .A2(_05406_),
    .ZN(_05439_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _11171_ (.A1(_02229_),
    .A2(_02261_),
    .A3(_04569_),
    .ZN(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11172_ (.I(_05440_),
    .Z(_05441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11173_ (.I(_05390_),
    .Z(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11174_ (.A1(net203),
    .A2(_05441_),
    .B(_05442_),
    .ZN(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11175_ (.A1(\as2650.chirpchar[1] ),
    .A2(_05377_),
    .ZN(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11176_ (.A1(_05439_),
    .A2(_05443_),
    .B(_05444_),
    .C(_05404_),
    .ZN(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11177_ (.A1(_05438_),
    .A2(_05445_),
    .ZN(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11178_ (.A1(_03007_),
    .A2(_05413_),
    .ZN(_05447_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11179_ (.A1(_05402_),
    .A2(_05446_),
    .B(_05447_),
    .C(_05434_),
    .ZN(_05448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11180_ (.A1(_02269_),
    .A2(_05435_),
    .B(_05448_),
    .ZN(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11181_ (.A1(_01860_),
    .A2(_05418_),
    .ZN(_05450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11182_ (.A1(_05399_),
    .A2(_05449_),
    .B(_05450_),
    .ZN(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11183_ (.A1(_05382_),
    .A2(_05451_),
    .B(_05388_),
    .ZN(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11184_ (.I(_05423_),
    .Z(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11185_ (.I(_05428_),
    .Z(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11186_ (.A1(_05347_),
    .A2(_05453_),
    .B1(_05454_),
    .B2(\as2650.regs[4][1] ),
    .ZN(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11187_ (.A1(_05433_),
    .A2(_05452_),
    .B(_05455_),
    .ZN(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11188_ (.I(_05387_),
    .Z(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11189_ (.A1(_01043_),
    .A2(_05432_),
    .ZN(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11190_ (.A1(_03086_),
    .A2(_05365_),
    .B(_05382_),
    .C(_05457_),
    .ZN(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11191_ (.I(_05398_),
    .Z(_05459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11192_ (.I(_05376_),
    .Z(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11193_ (.A1(net172),
    .A2(_05405_),
    .ZN(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11194_ (.A1(_04133_),
    .A2(_05407_),
    .B(_05461_),
    .C(_05391_),
    .ZN(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11195_ (.A1(\as2650.chirpchar[2] ),
    .A2(_05403_),
    .B(_05404_),
    .C(_05462_),
    .ZN(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11196_ (.A1(_05066_),
    .A2(_05411_),
    .ZN(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11197_ (.A1(_05463_),
    .A2(_05464_),
    .B(_05413_),
    .ZN(_05465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11198_ (.A1(_03069_),
    .A2(_05460_),
    .B(_05465_),
    .ZN(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11199_ (.A1(_02289_),
    .A2(_05416_),
    .ZN(_05467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11200_ (.I(_05398_),
    .Z(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11201_ (.A1(_05401_),
    .A2(_05466_),
    .B(_05467_),
    .C(_05468_),
    .ZN(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11202_ (.A1(_01869_),
    .A2(_05459_),
    .B(_05469_),
    .ZN(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11203_ (.A1(_05397_),
    .A2(_05470_),
    .ZN(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11204_ (.A1(_05456_),
    .A2(_05458_),
    .A3(_05471_),
    .ZN(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11205_ (.A1(_05349_),
    .A2(_05424_),
    .B1(_05429_),
    .B2(\as2650.regs[4][2] ),
    .ZN(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11206_ (.A1(_05472_),
    .A2(_05473_),
    .ZN(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11207_ (.I(_05381_),
    .Z(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11208_ (.A1(\as2650.regs[0][3] ),
    .A2(_05432_),
    .ZN(_05475_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11209_ (.A1(_03136_),
    .A2(_05365_),
    .B(_05474_),
    .C(_05475_),
    .ZN(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11210_ (.A1(_04188_),
    .A2(_05440_),
    .ZN(_05477_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11211_ (.A1(_02427_),
    .A2(_05440_),
    .B(_05477_),
    .C(_05390_),
    .ZN(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11212_ (.A1(\as2650.chirpchar[3] ),
    .A2(_05403_),
    .B(_05404_),
    .C(_05478_),
    .ZN(_05479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11213_ (.A1(_05065_),
    .A2(_05411_),
    .ZN(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11214_ (.A1(_05479_),
    .A2(_05480_),
    .B(_05413_),
    .ZN(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11215_ (.A1(_03117_),
    .A2(_05460_),
    .B(_05481_),
    .ZN(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11216_ (.A1(_01804_),
    .A2(_05400_),
    .ZN(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11217_ (.A1(_05416_),
    .A2(_05482_),
    .B(_05483_),
    .C(_05468_),
    .ZN(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11218_ (.A1(_01881_),
    .A2(_05459_),
    .B(_05484_),
    .ZN(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11219_ (.A1(_05397_),
    .A2(_05485_),
    .ZN(_05486_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11220_ (.A1(_05456_),
    .A2(_05476_),
    .A3(_05486_),
    .ZN(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11221_ (.A1(_05351_),
    .A2(_05424_),
    .B1(_05429_),
    .B2(\as2650.regs[4][3] ),
    .ZN(_05488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11222_ (.A1(_05487_),
    .A2(_05488_),
    .ZN(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11223_ (.I(_05378_),
    .Z(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11224_ (.A1(_05064_),
    .A2(_05489_),
    .ZN(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11225_ (.I(_05393_),
    .Z(_05491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11226_ (.I(_05405_),
    .Z(_05492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11227_ (.A1(net174),
    .A2(_05406_),
    .ZN(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11228_ (.A1(_04231_),
    .A2(_05492_),
    .B(_05493_),
    .C(_05442_),
    .ZN(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11229_ (.A1(\as2650.chirpchar[4] ),
    .A2(_05403_),
    .B(_05491_),
    .C(_05494_),
    .ZN(_05495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11230_ (.A1(_05490_),
    .A2(_05495_),
    .B(_05402_),
    .ZN(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _11231_ (.A1(_03176_),
    .A2(_05402_),
    .B(_05401_),
    .C(_05496_),
    .ZN(_05497_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11232_ (.A1(_01814_),
    .A2(_05435_),
    .B(_05418_),
    .ZN(_05498_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _11233_ (.A1(_05264_),
    .A2(_05399_),
    .B1(_05497_),
    .B2(_05498_),
    .ZN(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11234_ (.A1(\as2650.regs[0][4] ),
    .A2(_05367_),
    .ZN(_05500_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11235_ (.A1(_03187_),
    .A2(_05364_),
    .B(_05381_),
    .C(_05500_),
    .ZN(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11236_ (.A1(_05382_),
    .A2(_05499_),
    .B(_05501_),
    .C(_05388_),
    .ZN(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11237_ (.A1(_05354_),
    .A2(_05424_),
    .B1(_05429_),
    .B2(\as2650.regs[4][4] ),
    .ZN(_05503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11238_ (.A1(_05502_),
    .A2(_05503_),
    .ZN(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11239_ (.A1(\as2650.regs[0][5] ),
    .A2(_05367_),
    .ZN(_05504_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11240_ (.A1(_03232_),
    .A2(_05364_),
    .B(_05474_),
    .C(_05504_),
    .ZN(_05505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11241_ (.A1(\as2650.chirpchar[5] ),
    .A2(_05377_),
    .ZN(_05506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11242_ (.A1(_02451_),
    .A2(_05407_),
    .ZN(_05507_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11243_ (.A1(_04272_),
    .A2(_05406_),
    .B(_05507_),
    .C(_05391_),
    .ZN(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11244_ (.A1(_05506_),
    .A2(_05508_),
    .B(_05437_),
    .ZN(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _11245_ (.A1(_05062_),
    .A2(_05489_),
    .B(_05509_),
    .C(_05460_),
    .ZN(_05510_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11246_ (.A1(_03216_),
    .A2(_05389_),
    .B(_05434_),
    .ZN(_05511_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _11247_ (.A1(_01466_),
    .A2(_05435_),
    .B1(_05510_),
    .B2(_05511_),
    .C(_05468_),
    .ZN(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11248_ (.A1(_01897_),
    .A2(_05399_),
    .B(_05512_),
    .ZN(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11249_ (.A1(_05397_),
    .A2(_05513_),
    .ZN(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11250_ (.A1(_05456_),
    .A2(_05505_),
    .A3(_05514_),
    .ZN(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11251_ (.A1(_05358_),
    .A2(_05453_),
    .B1(_05454_),
    .B2(\as2650.regs[4][5] ),
    .ZN(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11252_ (.A1(_05515_),
    .A2(_05516_),
    .ZN(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11253_ (.A1(\as2650.regs[0][6] ),
    .A2(_05367_),
    .ZN(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11254_ (.A1(_03284_),
    .A2(_05364_),
    .B(_05474_),
    .C(_05517_),
    .ZN(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11255_ (.A1(_02460_),
    .A2(_05407_),
    .ZN(_05519_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11256_ (.A1(_04304_),
    .A2(_05492_),
    .B(_05519_),
    .C(_05442_),
    .ZN(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11257_ (.A1(\as2650.chirpchar[6] ),
    .A2(_05377_),
    .B(_05411_),
    .ZN(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11258_ (.A1(_05061_),
    .A2(_05437_),
    .B1(_05520_),
    .B2(_05521_),
    .C(_05376_),
    .ZN(_05522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11259_ (.A1(_03267_),
    .A2(_05460_),
    .B(_05522_),
    .ZN(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11260_ (.A1(_05401_),
    .A2(_05523_),
    .ZN(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11261_ (.A1(_04726_),
    .A2(_05435_),
    .B(_05418_),
    .ZN(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _11262_ (.A1(_01903_),
    .A2(_05459_),
    .B1(_05524_),
    .B2(_05525_),
    .ZN(_05526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11263_ (.A1(_05396_),
    .A2(_05526_),
    .ZN(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11264_ (.A1(_05388_),
    .A2(_05518_),
    .A3(_05527_),
    .ZN(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11265_ (.A1(_05360_),
    .A2(_05453_),
    .B1(_05454_),
    .B2(\as2650.regs[4][6] ),
    .ZN(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11266_ (.A1(_05528_),
    .A2(_05529_),
    .ZN(_00521_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11267_ (.A1(net177),
    .A2(_05441_),
    .B(_05393_),
    .C(_05442_),
    .ZN(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11268_ (.A1(_04349_),
    .A2(_05441_),
    .B(_05530_),
    .ZN(_05531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11269_ (.A1(_05060_),
    .A2(_05491_),
    .B(_05389_),
    .ZN(_05532_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _11270_ (.A1(_03329_),
    .A2(_05389_),
    .B1(_05531_),
    .B2(_05532_),
    .C(_05434_),
    .ZN(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11271_ (.A1(_01468_),
    .A2(_05416_),
    .ZN(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11272_ (.A1(_05468_),
    .A2(_05533_),
    .A3(_05534_),
    .ZN(_05535_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11273_ (.A1(_01910_),
    .A2(_05459_),
    .B(_05535_),
    .ZN(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11274_ (.A1(\as2650.regs[0][7] ),
    .A2(_05432_),
    .ZN(_05537_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11275_ (.A1(_03327_),
    .A2(_05365_),
    .B1(_05474_),
    .B2(_05536_),
    .C(_05537_),
    .ZN(_05538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11276_ (.A1(_05456_),
    .A2(_05538_),
    .ZN(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11277_ (.A1(_05362_),
    .A2(_05453_),
    .B1(_05454_),
    .B2(\as2650.regs[4][7] ),
    .ZN(_05540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11278_ (.A1(_05539_),
    .A2(_05540_),
    .ZN(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _11279_ (.A1(_01476_),
    .A2(_05334_),
    .ZN(_05541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11280_ (.A1(_00791_),
    .A2(_05541_),
    .ZN(_05542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11281_ (.I(_05542_),
    .Z(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11282_ (.I(_02947_),
    .Z(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _11283_ (.A1(_02825_),
    .A2(_05426_),
    .A3(_02963_),
    .ZN(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11284_ (.I(_05545_),
    .Z(_05546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11285_ (.I(_05393_),
    .Z(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11286_ (.I(_05547_),
    .Z(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11287_ (.I(_05440_),
    .Z(_05549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11288_ (.I(_05549_),
    .Z(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11289_ (.A1(_04387_),
    .A2(_05549_),
    .ZN(_05551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11290_ (.I(_05491_),
    .Z(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11291_ (.A1(net171),
    .A2(_05550_),
    .B(_05551_),
    .C(_05552_),
    .ZN(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11292_ (.A1(_05059_),
    .A2(_05548_),
    .B(_05553_),
    .ZN(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11293_ (.A1(_05491_),
    .A2(_05373_),
    .B(_02825_),
    .ZN(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11294_ (.I(_05555_),
    .Z(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11295_ (.I(_05542_),
    .ZN(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _11296_ (.A1(_02967_),
    .A2(_05557_),
    .A3(_05555_),
    .A4(_05545_),
    .ZN(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11297_ (.I(_05558_),
    .Z(_05559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11298_ (.A1(_05544_),
    .A2(_05546_),
    .B1(_05554_),
    .B2(_05556_),
    .C1(_05559_),
    .C2(\as2650.regs[1][0] ),
    .ZN(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11299_ (.A1(_02956_),
    .A2(_05543_),
    .B(_05560_),
    .ZN(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11300_ (.I(_05437_),
    .Z(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11301_ (.A1(_05058_),
    .A2(_05561_),
    .ZN(_05562_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11302_ (.I(_05441_),
    .Z(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11303_ (.A1(_04427_),
    .A2(_05563_),
    .ZN(_05564_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11304_ (.A1(net182),
    .A2(_05550_),
    .B(_05564_),
    .C(_05548_),
    .ZN(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11305_ (.A1(_05562_),
    .A2(_05565_),
    .ZN(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11306_ (.A1(_03037_),
    .A2(_05546_),
    .B1(_05566_),
    .B2(_05556_),
    .C1(_05559_),
    .C2(\as2650.regs[1][1] ),
    .ZN(_05567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11307_ (.A1(_03035_),
    .A2(_05543_),
    .B(_05567_),
    .ZN(_00524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11308_ (.I(_05545_),
    .Z(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11309_ (.I(_05558_),
    .Z(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11310_ (.A1(_05547_),
    .A2(_05373_),
    .ZN(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11311_ (.A1(_04665_),
    .A2(_05570_),
    .ZN(_05571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11312_ (.I(_05492_),
    .Z(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11313_ (.A1(net193),
    .A2(_05492_),
    .ZN(_05573_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11314_ (.A1(_04458_),
    .A2(_05572_),
    .B(_05573_),
    .C(_05547_),
    .ZN(_05574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11315_ (.A1(_05057_),
    .A2(_05548_),
    .B(_05574_),
    .ZN(_05575_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11316_ (.A1(_05571_),
    .A2(_05575_),
    .ZN(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11317_ (.A1(_03089_),
    .A2(_05568_),
    .B1(_05569_),
    .B2(\as2650.regs[1][2] ),
    .C(_05576_),
    .ZN(_05577_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11318_ (.A1(_03088_),
    .A2(_05543_),
    .B(_05577_),
    .ZN(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11319_ (.A1(_05056_),
    .A2(_05561_),
    .ZN(_05578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11320_ (.A1(_04493_),
    .A2(_05563_),
    .ZN(_05579_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11321_ (.A1(net197),
    .A2(_05550_),
    .B(_05579_),
    .C(_05548_),
    .ZN(_05580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11322_ (.A1(_05578_),
    .A2(_05580_),
    .ZN(_05581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11323_ (.A1(_03139_),
    .A2(_05546_),
    .B1(_05581_),
    .B2(_05556_),
    .C1(_05559_),
    .C2(\as2650.regs[1][3] ),
    .ZN(_05582_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11324_ (.A1(_03138_),
    .A2(_05543_),
    .B(_05582_),
    .ZN(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11325_ (.I(_05542_),
    .Z(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11326_ (.A1(_04529_),
    .A2(_05549_),
    .ZN(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11327_ (.A1(_02317_),
    .A2(_05563_),
    .B(_05584_),
    .C(_05552_),
    .ZN(_05585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11328_ (.A1(_05055_),
    .A2(_05561_),
    .ZN(_05586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11329_ (.A1(_05585_),
    .A2(_05586_),
    .ZN(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11330_ (.A1(_05571_),
    .A2(_05587_),
    .ZN(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11331_ (.A1(_03189_),
    .A2(_05568_),
    .B1(_05569_),
    .B2(\as2650.regs[1][4] ),
    .C(_05588_),
    .ZN(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11332_ (.A1(_03188_),
    .A2(_05583_),
    .B(_05589_),
    .ZN(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11333_ (.A1(net199),
    .A2(_05572_),
    .ZN(_05590_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11334_ (.A1(_03866_),
    .A2(_05572_),
    .B(_05590_),
    .C(_05552_),
    .ZN(_05591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11335_ (.A1(_05054_),
    .A2(_05489_),
    .ZN(_05592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11336_ (.A1(_05591_),
    .A2(_05592_),
    .ZN(_05593_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11337_ (.A1(_05571_),
    .A2(_05593_),
    .ZN(_05594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11338_ (.A1(_03234_),
    .A2(_05568_),
    .B1(_05569_),
    .B2(\as2650.regs[1][5] ),
    .C(_05594_),
    .ZN(_05595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11339_ (.A1(_03233_),
    .A2(_05583_),
    .B(_05595_),
    .ZN(_00528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11340_ (.A1(_03896_),
    .A2(_05549_),
    .ZN(_05596_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11341_ (.A1(_02346_),
    .A2(_05563_),
    .B(_05596_),
    .C(_05552_),
    .ZN(_05597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11342_ (.A1(_05053_),
    .A2(_05489_),
    .ZN(_05598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11343_ (.A1(_05597_),
    .A2(_05598_),
    .ZN(_05599_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11344_ (.A1(_05571_),
    .A2(_05599_),
    .ZN(_05600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11345_ (.A1(_03286_),
    .A2(_05568_),
    .B1(_05569_),
    .B2(\as2650.regs[1][6] ),
    .C(_05600_),
    .ZN(_05601_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11346_ (.A1(_03285_),
    .A2(_05583_),
    .B(_05601_),
    .ZN(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11347_ (.A1(net201),
    .A2(_05572_),
    .ZN(_05602_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11348_ (.A1(_03919_),
    .A2(_05550_),
    .B(_05561_),
    .ZN(_05603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _11349_ (.A1(_02484_),
    .A2(_05052_),
    .B1(_05602_),
    .B2(_05603_),
    .ZN(_05604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11350_ (.A1(_03330_),
    .A2(_05546_),
    .B1(_05604_),
    .B2(_05556_),
    .C1(_05559_),
    .C2(\as2650.regs[1][7] ),
    .ZN(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11351_ (.A1(_03328_),
    .A2(_05583_),
    .B(_05605_),
    .ZN(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11352_ (.A1(_04678_),
    .A2(_05541_),
    .ZN(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11353_ (.I(_05606_),
    .Z(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _11354_ (.A1(_05339_),
    .A2(_04609_),
    .A3(_02963_),
    .ZN(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11355_ (.I(_05608_),
    .Z(_05609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _11356_ (.A1(_04678_),
    .A2(_05541_),
    .B(_05608_),
    .C(_05343_),
    .ZN(_05610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11357_ (.I(_05610_),
    .Z(_05611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11358_ (.A1(_05544_),
    .A2(_05609_),
    .B1(_05611_),
    .B2(\as2650.regs[3][0] ),
    .ZN(_05612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11359_ (.A1(_02956_),
    .A2(_05607_),
    .B(_05612_),
    .ZN(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11360_ (.A1(_05347_),
    .A2(_05609_),
    .B1(_05611_),
    .B2(\as2650.regs[3][1] ),
    .ZN(_05613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11361_ (.A1(_03035_),
    .A2(_05607_),
    .B(_05613_),
    .ZN(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11362_ (.A1(_05349_),
    .A2(_05609_),
    .B1(_05611_),
    .B2(\as2650.regs[3][2] ),
    .ZN(_05614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11363_ (.A1(_03088_),
    .A2(_05607_),
    .B(_05614_),
    .ZN(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11364_ (.A1(_05351_),
    .A2(_05609_),
    .B1(_05611_),
    .B2(\as2650.regs[3][3] ),
    .ZN(_05615_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11365_ (.A1(_03138_),
    .A2(_05607_),
    .B(_05615_),
    .ZN(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11366_ (.I(_05606_),
    .Z(_05616_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11367_ (.I(_05608_),
    .Z(_05617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11368_ (.I(_05610_),
    .Z(_05618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11369_ (.A1(_05354_),
    .A2(_05617_),
    .B1(_05618_),
    .B2(\as2650.regs[3][4] ),
    .ZN(_05619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11370_ (.A1(_03188_),
    .A2(_05616_),
    .B(_05619_),
    .ZN(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11371_ (.A1(_05358_),
    .A2(_05617_),
    .B1(_05618_),
    .B2(\as2650.regs[3][5] ),
    .ZN(_05620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11372_ (.A1(_03233_),
    .A2(_05616_),
    .B(_05620_),
    .ZN(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11373_ (.A1(_05360_),
    .A2(_05617_),
    .B1(_05618_),
    .B2(\as2650.regs[3][6] ),
    .ZN(_05621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11374_ (.A1(_03285_),
    .A2(_05616_),
    .B(_05621_),
    .ZN(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11375_ (.A1(_05362_),
    .A2(_05617_),
    .B1(_05618_),
    .B2(\as2650.regs[3][7] ),
    .ZN(_05622_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11376_ (.A1(_03328_),
    .A2(_05616_),
    .B(_05622_),
    .ZN(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _11377_ (.A1(_02823_),
    .A2(_05335_),
    .A3(_05104_),
    .Z(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11378_ (.I(_05623_),
    .Z(_05624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11379_ (.A1(_05547_),
    .A2(_05373_),
    .B(_05425_),
    .ZN(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11380_ (.I(_05625_),
    .Z(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _11381_ (.A1(_05425_),
    .A2(_05426_),
    .A3(_02963_),
    .ZN(_05627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11382_ (.I(_05627_),
    .Z(_05628_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11383_ (.I(_05623_),
    .ZN(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _11384_ (.A1(_02967_),
    .A2(_05629_),
    .A3(_05625_),
    .A4(_05627_),
    .ZN(_05630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11385_ (.I(_05630_),
    .Z(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11386_ (.A1(_05554_),
    .A2(_05626_),
    .B1(_05628_),
    .B2(_05544_),
    .C1(\as2650.regs[5][0] ),
    .C2(_05631_),
    .ZN(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11387_ (.A1(_02955_),
    .A2(_05624_),
    .B(_05632_),
    .ZN(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11388_ (.A1(_05566_),
    .A2(_05626_),
    .B1(_05628_),
    .B2(_03037_),
    .C1(\as2650.regs[5][1] ),
    .C2(_05631_),
    .ZN(_05633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11389_ (.A1(_03034_),
    .A2(_05624_),
    .B(_05633_),
    .ZN(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11390_ (.I(_05627_),
    .Z(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11391_ (.I(_05630_),
    .Z(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11392_ (.A1(_01814_),
    .A2(_05570_),
    .ZN(_05636_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11393_ (.A1(_05575_),
    .A2(_05636_),
    .ZN(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11394_ (.A1(_03089_),
    .A2(_05634_),
    .B1(_05635_),
    .B2(\as2650.regs[5][2] ),
    .C(_05637_),
    .ZN(_05638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11395_ (.A1(_03087_),
    .A2(_05624_),
    .B(_05638_),
    .ZN(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11396_ (.A1(_05581_),
    .A2(_05626_),
    .B1(_05628_),
    .B2(_03139_),
    .C1(\as2650.regs[5][3] ),
    .C2(_05631_),
    .ZN(_05639_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11397_ (.A1(_03137_),
    .A2(_05624_),
    .B(_05639_),
    .ZN(_00542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11398_ (.I(_05623_),
    .Z(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11399_ (.A1(_05587_),
    .A2(_05636_),
    .ZN(_05641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11400_ (.A1(_03189_),
    .A2(_05634_),
    .B1(_05635_),
    .B2(\as2650.regs[5][4] ),
    .C(_05641_),
    .ZN(_05642_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11401_ (.A1(_03187_),
    .A2(_05640_),
    .B(_05642_),
    .ZN(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11402_ (.A1(_05593_),
    .A2(_05636_),
    .ZN(_05643_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11403_ (.A1(_03234_),
    .A2(_05634_),
    .B1(_05635_),
    .B2(\as2650.regs[5][5] ),
    .C(_05643_),
    .ZN(_05644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11404_ (.A1(_03232_),
    .A2(_05640_),
    .B(_05644_),
    .ZN(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11405_ (.A1(_05599_),
    .A2(_05636_),
    .ZN(_05645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11406_ (.A1(_03286_),
    .A2(_05634_),
    .B1(_05635_),
    .B2(\as2650.regs[5][6] ),
    .C(_05645_),
    .ZN(_05646_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11407_ (.A1(_03284_),
    .A2(_05640_),
    .B(_05646_),
    .ZN(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11408_ (.A1(_05604_),
    .A2(_05626_),
    .B1(_05628_),
    .B2(_03330_),
    .C1(\as2650.regs[5][7] ),
    .C2(_05631_),
    .ZN(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11409_ (.A1(_03327_),
    .A2(_05640_),
    .B(_05647_),
    .ZN(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11410_ (.A1(_02825_),
    .A2(_05426_),
    .A3(_05336_),
    .ZN(_05648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11411_ (.I(_05648_),
    .Z(_05649_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11412_ (.A1(_02964_),
    .A2(_05340_),
    .ZN(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11413_ (.I(_05650_),
    .Z(_05651_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11414_ (.I(_05648_),
    .ZN(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _11415_ (.A1(_05343_),
    .A2(_05650_),
    .A3(_05652_),
    .ZN(_05653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11416_ (.I(_05653_),
    .Z(_05654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11417_ (.A1(_05544_),
    .A2(_05651_),
    .B1(_05654_),
    .B2(\as2650.regs[6][0] ),
    .ZN(_05655_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11418_ (.A1(_02955_),
    .A2(_05649_),
    .B(_05655_),
    .ZN(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11419_ (.A1(_05347_),
    .A2(_05651_),
    .B1(_05654_),
    .B2(\as2650.regs[6][1] ),
    .ZN(_05656_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11420_ (.A1(_03034_),
    .A2(_05649_),
    .B(_05656_),
    .ZN(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11421_ (.A1(_03089_),
    .A2(_05651_),
    .B1(_05654_),
    .B2(\as2650.regs[6][2] ),
    .ZN(_05657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11422_ (.A1(_03087_),
    .A2(_05649_),
    .B(_05657_),
    .ZN(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11423_ (.A1(_03139_),
    .A2(_05651_),
    .B1(_05654_),
    .B2(\as2650.regs[6][3] ),
    .ZN(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11424_ (.A1(_03137_),
    .A2(_05649_),
    .B(_05658_),
    .ZN(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11425_ (.I(_05648_),
    .Z(_05659_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11426_ (.I(_05650_),
    .Z(_05660_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11427_ (.I(_05653_),
    .Z(_05661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11428_ (.A1(_03189_),
    .A2(_05660_),
    .B1(_05661_),
    .B2(\as2650.regs[6][4] ),
    .ZN(_05662_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11429_ (.A1(_03187_),
    .A2(_05659_),
    .B(_05662_),
    .ZN(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11430_ (.A1(_03234_),
    .A2(_05660_),
    .B1(_05661_),
    .B2(\as2650.regs[6][5] ),
    .ZN(_05663_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11431_ (.A1(_03232_),
    .A2(_05659_),
    .B(_05663_),
    .ZN(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11432_ (.A1(_03286_),
    .A2(_05660_),
    .B1(_05661_),
    .B2(\as2650.regs[6][6] ),
    .ZN(_05664_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11433_ (.A1(_03284_),
    .A2(_05659_),
    .B(_05664_),
    .ZN(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11434_ (.A1(_03330_),
    .A2(_05660_),
    .B1(_05661_),
    .B2(\as2650.regs[6][7] ),
    .ZN(_05665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11435_ (.A1(_03327_),
    .A2(_05659_),
    .B(_05665_),
    .ZN(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11436_ (.I(_05384_),
    .Z(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11437_ (.A1(_01618_),
    .A2(_05541_),
    .ZN(_05667_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11438_ (.I(_05667_),
    .Z(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11439_ (.A1(_05425_),
    .A2(_05380_),
    .ZN(_05669_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11440_ (.I(_05669_),
    .Z(_05670_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _11441_ (.A1(_00867_),
    .A2(_05666_),
    .B1(_05668_),
    .B2(_02954_),
    .C(_05670_),
    .ZN(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _11442_ (.A1(_04546_),
    .A2(_03677_),
    .A3(_05366_),
    .A4(_05385_),
    .ZN(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11443_ (.I(_05672_),
    .Z(_05673_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11444_ (.A1(_04665_),
    .A2(_05395_),
    .Z(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11445_ (.A1(_05420_),
    .A2(_05674_),
    .ZN(_05675_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11446_ (.A1(_05671_),
    .A2(_05673_),
    .A3(_05675_),
    .ZN(_05676_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _11447_ (.A1(_05339_),
    .A2(_02967_),
    .A3(_05386_),
    .ZN(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11448_ (.I(_05677_),
    .Z(_05678_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11449_ (.A1(_05366_),
    .A2(_05667_),
    .A3(_05669_),
    .A4(_05672_),
    .Z(_05679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11450_ (.I(_05679_),
    .Z(_05680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11451_ (.A1(_02957_),
    .A2(_05678_),
    .B1(_05680_),
    .B2(_01002_),
    .ZN(_05681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11452_ (.A1(_05676_),
    .A2(_05681_),
    .ZN(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _11453_ (.A1(_01478_),
    .A2(_01393_),
    .A3(_05335_),
    .ZN(_05682_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11454_ (.I(_05670_),
    .ZN(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11455_ (.A1(_00852_),
    .A2(_05666_),
    .ZN(_05684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11456_ (.A1(_05431_),
    .A2(_05682_),
    .B1(_05683_),
    .B2(_05451_),
    .C(_05684_),
    .ZN(_05685_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11457_ (.I(_05679_),
    .Z(_05686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11458_ (.A1(_03037_),
    .A2(_05677_),
    .B1(_05686_),
    .B2(_01020_),
    .ZN(_05687_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11459_ (.A1(_05678_),
    .A2(_05685_),
    .B(_05687_),
    .ZN(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11460_ (.I(_05673_),
    .Z(_05688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11461_ (.I(_05668_),
    .Z(_05689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11462_ (.I(_05669_),
    .Z(_05690_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11463_ (.A1(_04665_),
    .A2(_05343_),
    .ZN(_05691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11464_ (.A1(\as2650.regs[4][2] ),
    .A2(_05691_),
    .ZN(_05692_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _11465_ (.A1(_03087_),
    .A2(_05689_),
    .B1(_05690_),
    .B2(_05470_),
    .C(_05692_),
    .ZN(_05693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11466_ (.A1(_05688_),
    .A2(_05693_),
    .ZN(_05694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11467_ (.A1(_05349_),
    .A2(_05678_),
    .B1(_05680_),
    .B2(_01043_),
    .ZN(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11468_ (.A1(_05694_),
    .A2(_05695_),
    .ZN(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11469_ (.A1(\as2650.regs[4][3] ),
    .A2(_05691_),
    .ZN(_05696_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11470_ (.A1(_03137_),
    .A2(_05689_),
    .B1(_05690_),
    .B2(_05485_),
    .C(_05696_),
    .ZN(_05697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11471_ (.A1(_05688_),
    .A2(_05697_),
    .ZN(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11472_ (.A1(_05351_),
    .A2(_05678_),
    .B1(_05680_),
    .B2(\as2650.regs[0][3] ),
    .ZN(_05699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11473_ (.A1(_05698_),
    .A2(_05699_),
    .ZN(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11474_ (.A1(_00632_),
    .A2(_05666_),
    .B1(_05668_),
    .B2(_03186_),
    .C(_05669_),
    .ZN(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11475_ (.A1(_05499_),
    .A2(_05690_),
    .B(_05673_),
    .C(_05700_),
    .ZN(_05701_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11476_ (.I(_05677_),
    .Z(_05702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11477_ (.A1(_05354_),
    .A2(_05702_),
    .B1(_05680_),
    .B2(\as2650.regs[0][4] ),
    .ZN(_05703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11478_ (.A1(_05701_),
    .A2(_05703_),
    .ZN(_00559_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11479_ (.A1(_00816_),
    .A2(_05666_),
    .B1(_05668_),
    .B2(_03231_),
    .C(_05670_),
    .ZN(_05704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11480_ (.A1(_05513_),
    .A2(_05674_),
    .ZN(_05705_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11481_ (.A1(_05688_),
    .A2(_05704_),
    .A3(_05705_),
    .ZN(_05706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11482_ (.A1(_05358_),
    .A2(_05702_),
    .B1(_05686_),
    .B2(\as2650.regs[0][5] ),
    .ZN(_05707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11483_ (.A1(_05706_),
    .A2(_05707_),
    .ZN(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11484_ (.A1(\as2650.regs[4][6] ),
    .A2(_05691_),
    .ZN(_05708_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11485_ (.A1(_03283_),
    .A2(_05689_),
    .B(_05690_),
    .C(_05708_),
    .ZN(_05709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11486_ (.A1(_05526_),
    .A2(_05674_),
    .ZN(_05710_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11487_ (.A1(_05673_),
    .A2(_05709_),
    .A3(_05710_),
    .ZN(_05711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11488_ (.A1(_05360_),
    .A2(_05702_),
    .B1(_05686_),
    .B2(\as2650.regs[0][6] ),
    .ZN(_05712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11489_ (.A1(_05711_),
    .A2(_05712_),
    .ZN(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11490_ (.A1(\as2650.regs[4][7] ),
    .A2(_05691_),
    .ZN(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11491_ (.A1(_03326_),
    .A2(_05689_),
    .B1(_05670_),
    .B2(_05536_),
    .C(_05713_),
    .ZN(_05714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11492_ (.A1(_05688_),
    .A2(_05714_),
    .ZN(_05715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11493_ (.A1(_05362_),
    .A2(_05702_),
    .B1(_05686_),
    .B2(\as2650.regs[0][7] ),
    .ZN(_05716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11494_ (.A1(_05715_),
    .A2(_05716_),
    .ZN(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _11495_ (.A1(_02247_),
    .A2(_02248_),
    .A3(_02556_),
    .A4(_02599_),
    .ZN(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11496_ (.I(_05717_),
    .Z(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11497_ (.I0(_02555_),
    .I1(\as2650.stack[9][0] ),
    .S(_05718_),
    .Z(_05719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11498_ (.I(_05719_),
    .Z(_00563_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11499_ (.I0(_02560_),
    .I1(\as2650.stack[9][1] ),
    .S(_05718_),
    .Z(_05720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11500_ (.I(_05720_),
    .Z(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11501_ (.I0(_02562_),
    .I1(\as2650.stack[9][2] ),
    .S(_05718_),
    .Z(_05721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11502_ (.I(_05721_),
    .Z(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11503_ (.I0(_02564_),
    .I1(\as2650.stack[9][3] ),
    .S(_05718_),
    .Z(_05722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11504_ (.I(_05722_),
    .Z(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11505_ (.I(_05717_),
    .Z(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11506_ (.I0(_02566_),
    .I1(\as2650.stack[9][4] ),
    .S(_05723_),
    .Z(_05724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11507_ (.I(_05724_),
    .Z(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11508_ (.I0(_02569_),
    .I1(\as2650.stack[9][5] ),
    .S(_05723_),
    .Z(_05725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11509_ (.I(_05725_),
    .Z(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11510_ (.I0(_02571_),
    .I1(\as2650.stack[9][6] ),
    .S(_05723_),
    .Z(_05726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11511_ (.I(_05726_),
    .Z(_00569_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11512_ (.I0(_02573_),
    .I1(\as2650.stack[9][7] ),
    .S(_05723_),
    .Z(_05727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11513_ (.I(_05727_),
    .Z(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11514_ (.I(_05717_),
    .Z(_05728_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11515_ (.I0(_02575_),
    .I1(\as2650.stack[9][8] ),
    .S(_05728_),
    .Z(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11516_ (.I(_05729_),
    .Z(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11517_ (.I0(_02578_),
    .I1(\as2650.stack[9][9] ),
    .S(_05728_),
    .Z(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11518_ (.I(_05730_),
    .Z(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11519_ (.I0(_02580_),
    .I1(\as2650.stack[9][10] ),
    .S(_05728_),
    .Z(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11520_ (.I(_05731_),
    .Z(_00573_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11521_ (.I0(_02582_),
    .I1(\as2650.stack[9][11] ),
    .S(_05728_),
    .Z(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11522_ (.I(_05732_),
    .Z(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11523_ (.I(_05717_),
    .Z(_05733_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11524_ (.I0(_02584_),
    .I1(\as2650.stack[9][12] ),
    .S(_05733_),
    .Z(_05734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11525_ (.I(_05734_),
    .Z(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11526_ (.I0(_02587_),
    .I1(\as2650.stack[9][13] ),
    .S(_05733_),
    .Z(_05735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11527_ (.I(_05735_),
    .Z(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11528_ (.I0(_02589_),
    .I1(\as2650.stack[9][14] ),
    .S(_05733_),
    .Z(_05736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11529_ (.I(_05736_),
    .Z(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11530_ (.I0(_02591_),
    .I1(\as2650.stack[9][15] ),
    .S(_05733_),
    .Z(_05737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11531_ (.I(_05737_),
    .Z(_00578_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11532_ (.D(_00005_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.relative_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11533_ (.D(_00006_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(net106));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11534_ (.D(_00007_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(net113));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11535_ (.D(_00008_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(net114));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11536_ (.D(_00009_),
    .CLK(clknet_leaf_166_wb_clk_i),
    .Q(net115));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11537_ (.D(_00010_),
    .CLK(clknet_leaf_164_wb_clk_i),
    .Q(net116));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11538_ (.D(_00011_),
    .CLK(clknet_leaf_165_wb_clk_i),
    .Q(net117));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11539_ (.D(_00012_),
    .CLK(clknet_leaf_166_wb_clk_i),
    .Q(net118));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11540_ (.D(_00013_),
    .CLK(clknet_leaf_165_wb_clk_i),
    .Q(net119));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11541_ (.D(_00014_),
    .CLK(clknet_leaf_154_wb_clk_i),
    .Q(net120));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11542_ (.D(_00015_),
    .CLK(clknet_leaf_154_wb_clk_i),
    .Q(net121));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11543_ (.D(_00016_),
    .CLK(clknet_leaf_155_wb_clk_i),
    .Q(net107));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11544_ (.D(_00017_),
    .CLK(clknet_leaf_155_wb_clk_i),
    .Q(net108));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11545_ (.D(_00018_),
    .CLK(clknet_leaf_150_wb_clk_i),
    .Q(net109));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11546_ (.D(_00019_),
    .CLK(clknet_leaf_146_wb_clk_i),
    .Q(net110));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11547_ (.D(_00020_),
    .CLK(clknet_leaf_147_wb_clk_i),
    .Q(net111));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11548_ (.D(_00021_),
    .CLK(clknet_leaf_147_wb_clk_i),
    .Q(net112));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11549_ (.D(_00022_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(net90));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11550_ (.D(_00023_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(net97));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11551_ (.D(_00024_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(net98));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11552_ (.D(_00025_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(net99));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11553_ (.D(_00026_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(net100));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11554_ (.D(_00027_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(net101));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11555_ (.D(_00028_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(net102));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11556_ (.D(_00029_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(net103));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11557_ (.D(_00030_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(net104));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11558_ (.D(_00031_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(net105));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11559_ (.D(_00032_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(net91));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11560_ (.D(_00033_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(net92));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11561_ (.D(_00034_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(net93));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11562_ (.D(_00035_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(net94));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11563_ (.D(_00036_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(net95));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11564_ (.D(_00037_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(net96));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11565_ (.D(_00038_),
    .CLK(clknet_leaf_166_wb_clk_i),
    .Q(net142));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11566_ (.D(_00039_),
    .CLK(clknet_leaf_160_wb_clk_i),
    .Q(net143));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11567_ (.D(_00040_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(net144));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11568_ (.D(_00041_),
    .CLK(clknet_4_0__leaf_wb_clk_i),
    .Q(net215));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11569_ (.D(_00042_),
    .CLK(clknet_leaf_164_wb_clk_i),
    .Q(net216));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11570_ (.D(_00043_),
    .CLK(clknet_leaf_167_wb_clk_i),
    .Q(net227));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11571_ (.D(_00044_),
    .CLK(clknet_leaf_167_wb_clk_i),
    .Q(net238));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11572_ (.D(_00045_),
    .CLK(clknet_leaf_163_wb_clk_i),
    .Q(net241));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11573_ (.D(_00046_),
    .CLK(clknet_leaf_162_wb_clk_i),
    .Q(net242));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11574_ (.D(_00047_),
    .CLK(clknet_leaf_162_wb_clk_i),
    .Q(net243));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11575_ (.D(_00048_),
    .CLK(clknet_leaf_162_wb_clk_i),
    .Q(net244));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11576_ (.D(_00049_),
    .CLK(clknet_leaf_153_wb_clk_i),
    .Q(net245));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11577_ (.D(_00050_),
    .CLK(clknet_leaf_153_wb_clk_i),
    .Q(net246));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11578_ (.D(_00051_),
    .CLK(clknet_leaf_152_wb_clk_i),
    .Q(net247));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11579_ (.D(_00052_),
    .CLK(clknet_leaf_152_wb_clk_i),
    .Q(net217));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11580_ (.D(_00053_),
    .CLK(clknet_leaf_149_wb_clk_i),
    .Q(net218));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11581_ (.D(_00054_),
    .CLK(clknet_leaf_149_wb_clk_i),
    .Q(net219));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11582_ (.D(_00055_),
    .CLK(clknet_leaf_149_wb_clk_i),
    .Q(net220));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11583_ (.D(_00056_),
    .CLK(clknet_leaf_148_wb_clk_i),
    .Q(net221));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11584_ (.D(_00057_),
    .CLK(clknet_leaf_148_wb_clk_i),
    .Q(net222));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11585_ (.D(_00058_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(net223));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11586_ (.D(_00059_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(net224));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11587_ (.D(_00060_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(net225));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11588_ (.D(_00061_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(net226));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11589_ (.D(_00062_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(net228));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11590_ (.D(_00063_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(net229));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11591_ (.D(_00064_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(net230));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11592_ (.D(_00065_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(net231));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11593_ (.D(_00066_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(net232));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11594_ (.D(_00067_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(net233));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11595_ (.D(_00068_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(net234));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11596_ (.D(_00069_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(net235));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11597_ (.D(_00070_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(net236));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11598_ (.D(_00071_),
    .CLK(clknet_leaf_101_wb_clk_i),
    .Q(net237));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11599_ (.D(_00072_),
    .CLK(clknet_leaf_101_wb_clk_i),
    .Q(net239));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11600_ (.D(_00073_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(net240));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11601_ (.D(_00074_),
    .CLK(clknet_leaf_149_wb_clk_i),
    .Q(wb_feedback_delay));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11602_ (.D(net336),
    .CLK(clknet_leaf_159_wb_clk_i),
    .Q(wb_debug_cc));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11603_ (.D(net349),
    .CLK(clknet_leaf_159_wb_clk_i),
    .Q(wb_debug_carry));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11604_ (.D(net314),
    .CLK(clknet_leaf_160_wb_clk_i),
    .Q(\web_behavior[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11605_ (.D(net306),
    .CLK(clknet_leaf_160_wb_clk_i),
    .Q(\web_behavior[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11606_ (.D(net317),
    .CLK(clknet_leaf_161_wb_clk_i),
    .Q(wb_reset_override_en));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11607_ (.D(net324),
    .CLK(clknet_leaf_154_wb_clk_i),
    .Q(wb_reset_override));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11608_ (.D(_00081_),
    .CLK(clknet_leaf_160_wb_clk_i),
    .Q(wb_io3_test));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11609_ (.D(net320),
    .CLK(clknet_leaf_161_wb_clk_i),
    .Q(net165));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11610_ (.D(_00083_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\as2650.wb_hidden_rom_enable ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11611_ (.D(_00084_),
    .CLK(clknet_leaf_163_wb_clk_i),
    .Q(\wb_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11612_ (.D(_00085_),
    .CLK(clknet_leaf_163_wb_clk_i),
    .Q(\wb_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11613_ (.D(_00086_),
    .CLK(clknet_leaf_164_wb_clk_i),
    .Q(\wb_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11614_ (.D(_00087_),
    .CLK(clknet_leaf_163_wb_clk_i),
    .Q(\wb_counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11615_ (.D(_00088_),
    .CLK(clknet_leaf_161_wb_clk_i),
    .Q(\wb_counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11616_ (.D(_00089_),
    .CLK(clknet_leaf_161_wb_clk_i),
    .Q(\wb_counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11617_ (.D(_00090_),
    .CLK(clknet_leaf_162_wb_clk_i),
    .Q(\wb_counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11618_ (.D(_00091_),
    .CLK(clknet_leaf_153_wb_clk_i),
    .Q(\wb_counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11619_ (.D(net340),
    .CLK(clknet_leaf_154_wb_clk_i),
    .Q(\wb_counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11620_ (.D(net328),
    .CLK(clknet_leaf_152_wb_clk_i),
    .Q(\wb_counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11621_ (.D(net332),
    .CLK(clknet_leaf_152_wb_clk_i),
    .Q(\wb_counter[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11622_ (.D(net344),
    .CLK(clknet_leaf_150_wb_clk_i),
    .Q(\wb_counter[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11623_ (.D(net310),
    .CLK(clknet_leaf_149_wb_clk_i),
    .Q(\wb_counter[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11624_ (.D(_00097_),
    .CLK(clknet_leaf_148_wb_clk_i),
    .Q(\wb_counter[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11625_ (.D(_00098_),
    .CLK(clknet_leaf_148_wb_clk_i),
    .Q(\wb_counter[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11626_ (.D(_00099_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\wb_counter[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11627_ (.D(_00100_),
    .CLK(clknet_leaf_148_wb_clk_i),
    .Q(\wb_counter[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11628_ (.D(_00101_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\wb_counter[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11629_ (.D(_00102_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\wb_counter[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11630_ (.D(_00103_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\wb_counter[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11631_ (.D(_00104_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\wb_counter[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11632_ (.D(_00105_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\wb_counter[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11633_ (.D(_00106_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\wb_counter[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11634_ (.D(_00107_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\wb_counter[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11635_ (.D(_00108_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\wb_counter[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11636_ (.D(_00109_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\wb_counter[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11637_ (.D(_00110_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\wb_counter[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11638_ (.D(_00111_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(\wb_counter[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11639_ (.D(_00112_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(\wb_counter[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11640_ (.D(_00113_),
    .CLK(clknet_leaf_101_wb_clk_i),
    .Q(\wb_counter[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11641_ (.D(_00114_),
    .CLK(clknet_leaf_101_wb_clk_i),
    .Q(\wb_counter[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11642_ (.D(_00115_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\wb_counter[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11643_ (.D(_00116_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\as2650.chirpchar[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11644_ (.D(_00117_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.stack[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11645_ (.D(_00118_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\as2650.stack[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11646_ (.D(_00119_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.stack[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11647_ (.D(_00120_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11648_ (.D(_00121_),
    .CLK(clknet_leaf_157_wb_clk_i),
    .Q(\as2650.stack[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11649_ (.D(_00122_),
    .CLK(clknet_leaf_156_wb_clk_i),
    .Q(\as2650.stack[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11650_ (.D(_00123_),
    .CLK(clknet_leaf_157_wb_clk_i),
    .Q(\as2650.stack[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11651_ (.D(_00124_),
    .CLK(clknet_leaf_157_wb_clk_i),
    .Q(\as2650.stack[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11652_ (.D(_00125_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\as2650.stack[11][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11653_ (.D(_00126_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.stack[11][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11654_ (.D(_00127_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\as2650.stack[11][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11655_ (.D(_00128_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.stack[11][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11656_ (.D(_00129_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.stack[11][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11657_ (.D(_00130_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.stack[11][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11658_ (.D(_00131_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.stack[11][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11659_ (.D(_00132_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.stack[11][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11660_ (.D(_00133_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11661_ (.D(_00134_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11662_ (.D(_00135_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11663_ (.D(_00136_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11664_ (.D(_00137_),
    .CLK(clknet_leaf_159_wb_clk_i),
    .Q(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11665_ (.D(_00138_),
    .CLK(clknet_leaf_155_wb_clk_i),
    .Q(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11666_ (.D(_00139_),
    .CLK(clknet_leaf_156_wb_clk_i),
    .Q(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11667_ (.D(_00140_),
    .CLK(clknet_leaf_140_wb_clk_i),
    .Q(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11668_ (.D(_00141_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11669_ (.D(_00142_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11670_ (.D(_00143_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11671_ (.D(_00144_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11672_ (.D(_00145_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.stack[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11673_ (.D(_00146_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11674_ (.D(_00147_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.stack[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11675_ (.D(_00148_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[2][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11676_ (.D(_00149_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11677_ (.D(_00150_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11678_ (.D(_00151_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11679_ (.D(_00152_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11680_ (.D(_00153_),
    .CLK(clknet_leaf_158_wb_clk_i),
    .Q(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11681_ (.D(_00154_),
    .CLK(clknet_leaf_155_wb_clk_i),
    .Q(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11682_ (.D(_00155_),
    .CLK(clknet_leaf_156_wb_clk_i),
    .Q(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11683_ (.D(_00156_),
    .CLK(clknet_leaf_140_wb_clk_i),
    .Q(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11684_ (.D(_00157_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11685_ (.D(_00158_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11686_ (.D(_00159_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\as2650.stack[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11687_ (.D(_00160_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\as2650.stack[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11688_ (.D(_00161_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11689_ (.D(_00162_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11690_ (.D(_00163_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.stack[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11691_ (.D(_00164_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.stack[3][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11692_ (.D(_00165_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11693_ (.D(_00166_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11694_ (.D(_00167_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11695_ (.D(_00168_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11696_ (.D(_00169_),
    .CLK(clknet_leaf_159_wb_clk_i),
    .Q(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11697_ (.D(_00170_),
    .CLK(clknet_leaf_156_wb_clk_i),
    .Q(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11698_ (.D(_00171_),
    .CLK(clknet_leaf_156_wb_clk_i),
    .Q(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11699_ (.D(_00172_),
    .CLK(clknet_leaf_140_wb_clk_i),
    .Q(\as2650.stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11700_ (.D(_00173_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11701_ (.D(_00174_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11702_ (.D(_00175_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\as2650.stack[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11703_ (.D(_00176_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\as2650.stack[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11704_ (.D(_00177_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.stack[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11705_ (.D(_00178_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.stack[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11706_ (.D(_00179_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.stack[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11707_ (.D(_00180_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[0][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11708_ (.D(_00000_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\as2650.chirpchar[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11709_ (.D(_00001_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\as2650.chirpchar[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11710_ (.D(_00002_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\as2650.chirpchar[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11711_ (.D(_00003_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\as2650.chirpchar[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11712_ (.D(_00004_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\as2650.chirpchar[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11713_ (.D(_00181_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11714_ (.D(_00182_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11715_ (.D(_00183_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11716_ (.D(_00184_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11717_ (.D(_00185_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11718_ (.D(_00186_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11719_ (.D(_00187_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11720_ (.D(_00188_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11721_ (.D(_00189_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\as2650.stack[14][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11722_ (.D(_00190_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\as2650.stack[14][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11723_ (.D(_00191_),
    .CLK(clknet_leaf_136_wb_clk_i),
    .Q(\as2650.stack[14][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11724_ (.D(_00192_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(\as2650.stack[14][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11725_ (.D(_00193_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[14][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11726_ (.D(_00194_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.stack[14][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11727_ (.D(_00195_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.stack[14][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11728_ (.D(_00196_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[14][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11729_ (.D(_00197_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.stack[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11730_ (.D(_00198_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11731_ (.D(_00199_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.stack[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11732_ (.D(_00200_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\as2650.stack[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11733_ (.D(_00201_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11734_ (.D(_00202_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11735_ (.D(_00203_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11736_ (.D(_00204_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11737_ (.D(_00205_),
    .CLK(clknet_leaf_136_wb_clk_i),
    .Q(\as2650.stack[13][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11738_ (.D(_00206_),
    .CLK(clknet_leaf_135_wb_clk_i),
    .Q(\as2650.stack[13][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11739_ (.D(_00207_),
    .CLK(clknet_leaf_136_wb_clk_i),
    .Q(\as2650.stack[13][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11740_ (.D(_00208_),
    .CLK(clknet_leaf_135_wb_clk_i),
    .Q(\as2650.stack[13][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11741_ (.D(_00209_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[13][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11742_ (.D(_00210_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.stack[13][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11743_ (.D(_00211_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[13][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11744_ (.D(_00212_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.stack[13][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11745_ (.D(_00213_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(\as2650.stack[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11746_ (.D(_00214_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\as2650.stack[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11747_ (.D(_00215_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11748_ (.D(_00216_),
    .CLK(clknet_leaf_147_wb_clk_i),
    .Q(\as2650.stack[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11749_ (.D(_00217_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11750_ (.D(_00218_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11751_ (.D(_00219_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11752_ (.D(_00220_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11753_ (.D(_00221_),
    .CLK(clknet_leaf_136_wb_clk_i),
    .Q(\as2650.stack[12][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11754_ (.D(_00222_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(\as2650.stack[12][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11755_ (.D(_00223_),
    .CLK(clknet_leaf_139_wb_clk_i),
    .Q(\as2650.stack[12][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11756_ (.D(_00224_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(\as2650.stack[12][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11757_ (.D(_00225_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[12][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11758_ (.D(_00226_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.stack[12][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11759_ (.D(_00227_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.stack[12][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11760_ (.D(_00228_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.stack[12][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11761_ (.D(_00229_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(\as2650.stack[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11762_ (.D(_00230_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\as2650.stack[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11763_ (.D(_00231_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11764_ (.D(_00232_),
    .CLK(clknet_leaf_145_wb_clk_i),
    .Q(\as2650.stack[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11765_ (.D(_00233_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11766_ (.D(_00234_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11767_ (.D(_00235_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11768_ (.D(_00236_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11769_ (.D(_00237_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(\as2650.stack[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11770_ (.D(_00238_),
    .CLK(clknet_leaf_131_wb_clk_i),
    .Q(\as2650.stack[8][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11771_ (.D(_00239_),
    .CLK(clknet_4_3__leaf_wb_clk_i),
    .Q(\as2650.stack[8][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11772_ (.D(_00240_),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(\as2650.stack[8][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11773_ (.D(_00241_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[8][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11774_ (.D(_00242_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.stack[8][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11775_ (.D(_00243_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.stack[8][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11776_ (.D(_00244_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[8][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11777_ (.D(_00245_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11778_ (.D(_00246_),
    .CLK(clknet_leaf_142_wb_clk_i),
    .Q(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11779_ (.D(_00247_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11780_ (.D(_00248_),
    .CLK(clknet_leaf_145_wb_clk_i),
    .Q(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11781_ (.D(_00249_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11782_ (.D(_00250_),
    .CLK(clknet_leaf_160_wb_clk_i),
    .Q(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11783_ (.D(_00251_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11784_ (.D(_00252_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11785_ (.D(_00253_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.stack[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11786_ (.D(_00254_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.stack[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11787_ (.D(_00255_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.stack[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11788_ (.D(_00256_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.stack[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11789_ (.D(_00257_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.stack[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11790_ (.D(_00258_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11791_ (.D(_00259_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.stack[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11792_ (.D(_00260_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.stack[7][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11793_ (.D(_00261_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11794_ (.D(_00262_),
    .CLK(clknet_leaf_146_wb_clk_i),
    .Q(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11795_ (.D(_00263_),
    .CLK(clknet_leaf_142_wb_clk_i),
    .Q(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11796_ (.D(_00264_),
    .CLK(clknet_leaf_146_wb_clk_i),
    .Q(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11797_ (.D(_00265_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11798_ (.D(_00266_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11799_ (.D(_00267_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11800_ (.D(_00268_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11801_ (.D(_00269_),
    .CLK(clknet_leaf_139_wb_clk_i),
    .Q(\as2650.stack[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11802_ (.D(_00270_),
    .CLK(clknet_leaf_138_wb_clk_i),
    .Q(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11803_ (.D(_00271_),
    .CLK(clknet_leaf_138_wb_clk_i),
    .Q(\as2650.stack[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11804_ (.D(_00272_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.stack[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11805_ (.D(_00273_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11806_ (.D(_00274_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.stack[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11807_ (.D(_00275_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11808_ (.D(_00276_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.stack[6][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11809_ (.D(_00277_),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11810_ (.D(_00278_),
    .CLK(clknet_leaf_142_wb_clk_i),
    .Q(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11811_ (.D(_00279_),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11812_ (.D(_00280_),
    .CLK(clknet_leaf_155_wb_clk_i),
    .Q(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11813_ (.D(_00281_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11814_ (.D(_00282_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11815_ (.D(_00283_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11816_ (.D(_00284_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11817_ (.D(_00285_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11818_ (.D(_00286_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.stack[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11819_ (.D(_00287_),
    .CLK(clknet_leaf_138_wb_clk_i),
    .Q(\as2650.stack[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11820_ (.D(_00288_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.stack[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11821_ (.D(_00289_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11822_ (.D(_00290_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11823_ (.D(_00291_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11824_ (.D(_00292_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.stack[5][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11825_ (.D(_00293_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(\as2650.stack[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11826_ (.D(_00294_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11827_ (.D(_00295_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11828_ (.D(_00296_),
    .CLK(clknet_leaf_145_wb_clk_i),
    .Q(\as2650.stack[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11829_ (.D(_00297_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11830_ (.D(_00298_),
    .CLK(clknet_leaf_158_wb_clk_i),
    .Q(\as2650.stack[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11831_ (.D(_00299_),
    .CLK(clknet_leaf_157_wb_clk_i),
    .Q(\as2650.stack[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11832_ (.D(_00300_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11833_ (.D(_00301_),
    .CLK(clknet_leaf_131_wb_clk_i),
    .Q(\as2650.stack[10][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11834_ (.D(_00302_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\as2650.stack[10][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11835_ (.D(_00303_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(\as2650.stack[10][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11836_ (.D(_00304_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\as2650.stack[10][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11837_ (.D(_00305_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[10][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11838_ (.D(_00306_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[10][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11839_ (.D(_00307_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.stack[10][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11840_ (.D(_00308_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.stack[10][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11841_ (.D(_00309_),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11842_ (.D(_00310_),
    .CLK(clknet_4_2__leaf_wb_clk_i),
    .Q(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11843_ (.D(_00311_),
    .CLK(clknet_leaf_142_wb_clk_i),
    .Q(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11844_ (.D(_00312_),
    .CLK(clknet_leaf_155_wb_clk_i),
    .Q(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11845_ (.D(_00313_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11846_ (.D(_00314_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11847_ (.D(_00315_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11848_ (.D(_00316_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11849_ (.D(_00317_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11850_ (.D(_00318_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11851_ (.D(_00319_),
    .CLK(clknet_leaf_139_wb_clk_i),
    .Q(\as2650.stack[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11852_ (.D(_00320_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.stack[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11853_ (.D(_00321_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11854_ (.D(_00322_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.stack[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11855_ (.D(_00323_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.stack[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11856_ (.D(_00324_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.stack[4][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11857_ (.D(_00325_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(\as2650.stack[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11858_ (.D(_00326_),
    .CLK(clknet_leaf_145_wb_clk_i),
    .Q(\as2650.stack[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11859_ (.D(_00327_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(\as2650.stack[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11860_ (.D(_00328_),
    .CLK(clknet_leaf_145_wb_clk_i),
    .Q(\as2650.stack[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11861_ (.D(_00329_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11862_ (.D(_00330_),
    .CLK(clknet_leaf_158_wb_clk_i),
    .Q(\as2650.stack[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11863_ (.D(_00331_),
    .CLK(clknet_leaf_158_wb_clk_i),
    .Q(\as2650.stack[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11864_ (.D(_00332_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11865_ (.D(_00333_),
    .CLK(clknet_leaf_135_wb_clk_i),
    .Q(\as2650.stack[15][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11866_ (.D(_00334_),
    .CLK(clknet_leaf_135_wb_clk_i),
    .Q(\as2650.stack[15][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11867_ (.D(_00335_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(\as2650.stack[15][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11868_ (.D(_00336_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[15][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11869_ (.D(_00337_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[15][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11870_ (.D(_00338_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.stack[15][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11871_ (.D(_00339_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.stack[15][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11872_ (.D(_00340_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.stack[15][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11873_ (.D(_00341_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.regs[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11874_ (.D(_00342_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.regs[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11875_ (.D(_00343_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.regs[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11876_ (.D(_00344_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.regs[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11877_ (.D(_00345_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.regs[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11878_ (.D(_00346_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\as2650.regs[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11879_ (.D(_00347_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\as2650.regs[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11880_ (.D(_00348_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.regs[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11881_ (.D(_00349_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11882_ (.D(_00350_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11883_ (.D(_00351_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.stack[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11884_ (.D(_00352_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11885_ (.D(_00353_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11886_ (.D(_00354_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11887_ (.D(_00355_),
    .CLK(clknet_leaf_160_wb_clk_i),
    .Q(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11888_ (.D(_00356_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11889_ (.D(_00357_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\as2650.stack[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11890_ (.D(_00358_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\as2650.stack[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11891_ (.D(_00359_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\as2650.stack[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11892_ (.D(_00360_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\as2650.stack[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11893_ (.D(_00361_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11894_ (.D(_00362_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11895_ (.D(_00363_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.stack[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11896_ (.D(_00364_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[1][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11897_ (.D(_00365_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.last_addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11898_ (.D(_00366_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.last_addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11899_ (.D(_00367_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.last_addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11900_ (.D(_00368_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.last_addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11901_ (.D(_00369_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.last_addr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11902_ (.D(_00370_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.last_addr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11903_ (.D(_00371_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.last_addr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11904_ (.D(_00372_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.last_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11905_ (.D(_00373_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\as2650.chirp_ptr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11906_ (.D(_00374_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.chirp_ptr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11907_ (.D(_00375_),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(\as2650.chirp_ptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11908_ (.D(_00376_),
    .CLK(clknet_4_7__leaf_wb_clk_i),
    .Q(\as2650.indirect_target[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11909_ (.D(_00377_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.indirect_target[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11910_ (.D(_00378_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.indirect_target[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11911_ (.D(_00379_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.indirect_target[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11912_ (.D(_00380_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.indirect_target[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11913_ (.D(_00381_),
    .CLK(clknet_4_5__leaf_wb_clk_i),
    .Q(\as2650.indirect_target[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11914_ (.D(_00382_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.indirect_target[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11915_ (.D(_00383_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.indirect_target[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11916_ (.D(_00384_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.indirect_target[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11917_ (.D(_00385_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.indirect_target[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11918_ (.D(_00386_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.indirect_target[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11919_ (.D(_00387_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.indirect_target[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11920_ (.D(_00388_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.indirect_target[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11921_ (.D(_00389_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.indirect_target[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11922_ (.D(_00390_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.indirect_target[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11923_ (.D(_00391_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.indirect_target[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11924_ (.D(_00392_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.indexed_cyc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11925_ (.D(_00393_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.indexed_cyc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11926_ (.D(_00394_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.indirect_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11927_ (.D(_00395_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(net196));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11928_ (.D(_00396_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.extend ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11929_ (.D(_00397_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.warmup[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11930_ (.D(_00398_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.warmup[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11931_ (.D(_00399_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.instruction_args_latch[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11932_ (.D(_00400_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.instruction_args_latch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11933_ (.D(_00401_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.instruction_args_latch[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11934_ (.D(_00402_),
    .CLK(clknet_4_7__leaf_wb_clk_i),
    .Q(\as2650.instruction_args_latch[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11935_ (.D(_00403_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.instruction_args_latch[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11936_ (.D(_00404_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.instruction_args_latch[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11937_ (.D(_00405_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.instruction_args_latch[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11938_ (.D(_00406_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.instruction_args_latch[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11939_ (.D(_00407_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.instruction_args_latch[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11940_ (.D(_00408_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.instruction_args_latch[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11941_ (.D(_00409_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.instruction_args_latch[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11942_ (.D(_00410_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.instruction_args_latch[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11943_ (.D(_00411_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.instruction_args_latch[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11944_ (.D(_00412_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.instruction_args_latch[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11945_ (.D(_00413_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.instruction_args_latch[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11946_ (.D(_00414_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.instruction_args_latch[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11947_ (.D(_00415_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11948_ (.D(_00416_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11949_ (.D(_00417_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11950_ (.D(_00418_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11951_ (.D(_00419_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.insin[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11952_ (.D(_00420_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.insin[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11953_ (.D(_00421_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.insin[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11954_ (.D(_00422_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.insin[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11955_ (.D(_00423_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\as2650.insin[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11956_ (.D(_00424_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.insin[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11957_ (.D(_00425_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.insin[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11958_ (.D(_00426_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\as2650.insin[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11959_ (.D(_00427_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.page_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11960_ (.D(_00428_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.page_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11961_ (.D(_00429_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.page_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11962_ (.D(_00430_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.last_addr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11963_ (.D(_00431_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.last_addr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11964_ (.D(_00432_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.last_addr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11965_ (.D(_00433_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.last_addr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11966_ (.D(_00434_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.last_addr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11967_ (.D(_00435_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.last_addr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11968_ (.D(_00436_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.last_addr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11969_ (.D(_00437_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.last_addr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11970_ (.D(_00438_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.ivectors_base[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11971_ (.D(_00439_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.ivectors_base[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11972_ (.D(_00440_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.ivectors_base[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11973_ (.D(_00441_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.ivectors_base[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11974_ (.D(_00442_),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(\as2650.ivectors_base[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11975_ (.D(_00443_),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(\as2650.ivectors_base[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11976_ (.D(_00444_),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(\as2650.ivectors_base[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11977_ (.D(_00445_),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(\as2650.ivectors_base[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11978_ (.D(_00446_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.ivectors_base[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11979_ (.D(_00447_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.ivectors_base[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11980_ (.D(_00448_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.ivectors_base[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11981_ (.D(_00449_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.ivectors_base[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11982_ (.D(_00450_),
    .CLK(clknet_4_6__leaf_wb_clk_i),
    .Q(\as2650.PC[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11983_ (.D(_00451_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.PC[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11984_ (.D(_00452_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.PC[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11985_ (.D(_00453_),
    .CLK(clknet_4_6__leaf_wb_clk_i),
    .Q(\as2650.PC[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11986_ (.D(_00454_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.PC[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11987_ (.D(_00455_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.PC[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11988_ (.D(_00456_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.PC[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11989_ (.D(_00457_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.PC[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11990_ (.D(_00458_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.PC[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11991_ (.D(_00459_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.PC[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11992_ (.D(_00460_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.PC[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11993_ (.D(_00461_),
    .CLK(clknet_4_4__leaf_wb_clk_i),
    .Q(\as2650.PC[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11994_ (.D(_00462_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.PC[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11995_ (.D(_00463_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\as2650.debug_psl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11996_ (.D(_00464_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\as2650.debug_psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11997_ (.D(_00465_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.debug_psl[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11998_ (.D(_00466_),
    .CLK(clknet_4_12__leaf_wb_clk_i),
    .Q(\as2650.debug_psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11999_ (.D(_00467_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\as2650.debug_psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12000_ (.D(_00468_),
    .CLK(clknet_4_13__leaf_wb_clk_i),
    .Q(\as2650.debug_psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12001_ (.D(_00469_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\as2650.debug_psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12002_ (.D(_00470_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\as2650.debug_psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12003_ (.D(_00471_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.debug_psu[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12004_ (.D(_00472_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.debug_psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12005_ (.D(_00473_),
    .CLK(clknet_4_6__leaf_wb_clk_i),
    .Q(\as2650.debug_psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12006_ (.D(_00474_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.debug_psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12007_ (.D(_00475_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.debug_psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12008_ (.D(_00476_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.debug_psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12009_ (.D(_00477_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(net164));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12010_ (.D(_00478_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.debug_psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12011_ (.D(_00479_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.irqs_latch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12012_ (.D(_00480_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.irqs_latch[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12013_ (.D(_00481_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.irqs_latch[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12014_ (.D(_00482_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.irqs_latch[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12015_ (.D(_00483_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.irqs_latch[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12016_ (.D(_00484_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.irqs_latch[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12017_ (.D(_00485_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.irqs_latch[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12018_ (.D(_00486_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.trap ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12019_ (.D(_00487_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(net131));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12020_ (.D(_00488_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(net132));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12021_ (.D(_00489_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(net133));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12022_ (.D(_00490_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(net134));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12023_ (.D(_00491_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(net135));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12024_ (.D(_00492_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(net136));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12025_ (.D(_00493_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(net137));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12026_ (.D(_00494_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(net138));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12027_ (.D(_00495_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(net130));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12028_ (.D(_00496_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(net124));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12029_ (.D(_00497_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(net125));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12030_ (.D(_00498_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(net126));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12031_ (.D(_00499_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(net127));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12032_ (.D(_00500_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(net128));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12033_ (.D(_00501_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(net129));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12034_ (.D(_00502_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.ext_io_addr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12035_ (.D(_00503_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.ext_io_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12036_ (.D(_00504_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.io_bus_we ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12037_ (.D(_00505_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\as2650.chirpchar[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12038_ (.D(_00506_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.cpu_hidden_rom_enable ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12039_ (.D(_00507_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.regs[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12040_ (.D(_00508_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\as2650.regs[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12041_ (.D(_00509_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\as2650.regs[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12042_ (.D(_00510_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\as2650.regs[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12043_ (.D(_00511_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.regs[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12044_ (.D(_00512_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.regs[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12045_ (.D(_00513_),
    .CLK(clknet_4_14__leaf_wb_clk_i),
    .Q(\as2650.regs[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12046_ (.D(_00514_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\as2650.regs[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12047_ (.D(_00515_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\as2650.regs[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12048_ (.D(_00516_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.regs[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12049_ (.D(_00517_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\as2650.regs[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12050_ (.D(_00518_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\as2650.regs[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12051_ (.D(_00519_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(\as2650.regs[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12052_ (.D(_00520_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\as2650.regs[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12053_ (.D(_00521_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(\as2650.regs[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12054_ (.D(_00522_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12055_ (.D(_00523_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.regs[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12056_ (.D(_00524_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.regs[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12057_ (.D(_00525_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.regs[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12058_ (.D(_00526_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.regs[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12059_ (.D(_00527_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\as2650.regs[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12060_ (.D(_00528_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.regs[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12061_ (.D(_00529_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\as2650.regs[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12062_ (.D(_00530_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\as2650.regs[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12063_ (.D(_00531_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\as2650.regs[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12064_ (.D(_00532_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\as2650.regs[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12065_ (.D(_00533_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\as2650.regs[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12066_ (.D(_00534_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.regs[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12067_ (.D(_00535_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.regs[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12068_ (.D(_00536_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.regs[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12069_ (.D(_00537_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.regs[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12070_ (.D(_00538_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.regs[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12071_ (.D(_00539_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.regs[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12072_ (.D(_00540_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12073_ (.D(_00541_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\as2650.regs[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12074_ (.D(_00542_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\as2650.regs[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12075_ (.D(_00543_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.regs[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12076_ (.D(_00544_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.regs[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12077_ (.D(_00545_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.regs[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12078_ (.D(_00546_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.regs[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12079_ (.D(_00547_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\as2650.regs[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12080_ (.D(_00548_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\as2650.regs[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12081_ (.D(_00549_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\as2650.regs[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12082_ (.D(_00550_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\as2650.regs[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12083_ (.D(_00551_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\as2650.regs[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12084_ (.D(_00552_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\as2650.regs[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12085_ (.D(_00553_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\as2650.regs[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12086_ (.D(_00554_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\as2650.regs[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12087_ (.D(_00555_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\as2650.regs[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12088_ (.D(_00556_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.regs[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12089_ (.D(_00557_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\as2650.regs[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12090_ (.D(_00558_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\as2650.regs[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12091_ (.D(_00559_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(\as2650.regs[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12092_ (.D(_00560_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12093_ (.D(_00561_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(\as2650.regs[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12094_ (.D(_00562_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.regs[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12095_ (.D(_00563_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12096_ (.D(_00564_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12097_ (.D(_00565_),
    .CLK(clknet_4_9__leaf_wb_clk_i),
    .Q(\as2650.stack[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12098_ (.D(_00566_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12099_ (.D(_00567_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12100_ (.D(_00568_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.stack[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12101_ (.D(_00569_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12102_ (.D(_00570_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12103_ (.D(_00571_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\as2650.stack[9][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12104_ (.D(_00572_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\as2650.stack[9][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12105_ (.D(_00573_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\as2650.stack[9][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12106_ (.D(_00574_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\as2650.stack[9][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12107_ (.D(_00575_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[9][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12108_ (.D(_00576_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.stack[9][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12109_ (.D(_00577_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[9][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12110_ (.D(_00578_),
    .CLK(clknet_4_4__leaf_wb_clk_i),
    .Q(\as2650.stack[9][15] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12149_ (.I(net249),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12150_ (.I(net249),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12151_ (.I(net249),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12152_ (.I(net250),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12153_ (.I(net250),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12154_ (.I(net250),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12155_ (.I(net251),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12156_ (.I(net249),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12157_ (.I(net166),
    .Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12158_ (.I(net167),
    .Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12159_ (.I(net168),
    .Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12160_ (.I(net169),
    .Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12161_ (.I(net170),
    .Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12162_ (.I(net154),
    .Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12163_ (.I(net155),
    .Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12164_ (.I(net156),
    .Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_0__f_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_10__f_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_11__f_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_12__f_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_13__f_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_14__f_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_15__f_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_1__f_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_2__f_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_3__f_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_4__f_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_5__f_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_6__f_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_7__f_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_8__f_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_9__f_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_101_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_101_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_102_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_102_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_103_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_103_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_104_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_104_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_105_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_105_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_106_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_106_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_107_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_107_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_108_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_108_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_109_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_109_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_10_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_110_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_110_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_111_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_111_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_112_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_112_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_113_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_113_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_114_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_114_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_115_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_115_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_116_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_116_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_117_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_117_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_118_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_118_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_119_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_119_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_120_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_120_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_121_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_121_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_122_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_122_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_123_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_123_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_124_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_124_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_125_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_125_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_126_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_126_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_127_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_127_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_128_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_128_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_130_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_130_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_131_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_131_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_132_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_132_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_133_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_133_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_134_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_134_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_135_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_135_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_136_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_136_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_137_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_137_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_138_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_138_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_139_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_139_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_140_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_140_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_141_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_141_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_142_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_142_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_143_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_143_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_144_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_144_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_145_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_145_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_146_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_146_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_147_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_147_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_148_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_148_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_149_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_149_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_150_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_150_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_152_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_152_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_153_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_153_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_154_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_154_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_155_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_155_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_156_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_156_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_157_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_157_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_158_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_158_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_159_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_159_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_160_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_160_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_161_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_161_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_162_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_162_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_163_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_163_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_164_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_164_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_165_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_165_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_166_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_166_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_167_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_167_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_16_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_19_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_22_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_72_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_75_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_78_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_79_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_79_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_80_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_81_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_81_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_82_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_82_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_83_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_83_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_85_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_85_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_87_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_87_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_88_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_88_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_89_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_89_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_8_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_90_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_90_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_91_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_91_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_92_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_92_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_93_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_93_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_94_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_94_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_95_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_95_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_96_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_96_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_97_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_97_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_98_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_98_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_99_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_99_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout249 (.I(net250),
    .Z(net249));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout250 (.I(net147),
    .Z(net250));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout251 (.I(net147),
    .Z(net251));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 fanout253 (.I(net164),
    .Z(net253));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold100 (.I(wbs_dat_i[17]),
    .Z(net394));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold101 (.I(wbs_dat_i[7]),
    .Z(net395));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold102 (.I(wbs_dat_i[20]),
    .Z(net396));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold103 (.I(wbs_dat_i[2]),
    .Z(net397));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold104 (.I(wbs_dat_i[0]),
    .Z(net398));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold105 (.I(wbs_dat_i[22]),
    .Z(net399));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold106 (.I(wbs_dat_i[9]),
    .Z(net400));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold107 (.I(wbs_dat_i[21]),
    .Z(net401));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold108 (.I(wbs_dat_i[24]),
    .Z(net402));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold109 (.I(wbs_dat_i[23]),
    .Z(net403));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold11 (.I(net406),
    .Z(net303));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold110 (.I(wbs_dat_i[27]),
    .Z(net404));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold111 (.I(wbs_dat_i[25]),
    .Z(net405));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold112 (.I(wbs_dat_i[3]),
    .Z(net406));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold113 (.I(wbs_dat_i[26]),
    .Z(net407));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold114 (.I(wbs_dat_i[30]),
    .Z(net408));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold115 (.I(wbs_dat_i[1]),
    .Z(net409));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold116 (.I(wbs_dat_i[5]),
    .Z(net410));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold117 (.I(wbs_dat_i[28]),
    .Z(net411));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold118 (.I(wbs_dat_i[31]),
    .Z(net412));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold119 (.I(wbs_dat_i[18]),
    .Z(net413));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold12 (.I(net81),
    .Z(net304));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold120 (.I(wbs_adr_i[19]),
    .Z(net414));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold13 (.I(_02000_),
    .Z(net305));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold14 (.I(_00078_),
    .Z(net306));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold15 (.I(net359),
    .Z(net307));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold16 (.I(net59),
    .Z(net308));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold17 (.I(_02066_),
    .Z(net309));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold18 (.I(_00096_),
    .Z(net310));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold19 (.I(net397),
    .Z(net311));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold20 (.I(net78),
    .Z(net312));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold21 (.I(_01998_),
    .Z(net313));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold22 (.I(_00077_),
    .Z(net314));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold23 (.I(net382),
    .Z(net315));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold24 (.I(_02003_),
    .Z(net316));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold25 (.I(_00079_),
    .Z(net317));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold26 (.I(net395),
    .Z(net318));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold27 (.I(_02008_),
    .Z(net319));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold28 (.I(_00082_),
    .Z(net320));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold29 (.I(net410),
    .Z(net321));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold30 (.I(net83),
    .Z(net322));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold31 (.I(_02005_),
    .Z(net323));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold32 (.I(_00080_),
    .Z(net324));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold33 (.I(net400),
    .Z(net325));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold34 (.I(net87),
    .Z(net326));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold35 (.I(_02052_),
    .Z(net327));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold36 (.I(_00093_),
    .Z(net328));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold37 (.I(net383),
    .Z(net329));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold38 (.I(net57),
    .Z(net330));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold39 (.I(_02055_),
    .Z(net331));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold40 (.I(_00094_),
    .Z(net332));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold41 (.I(net398),
    .Z(net333));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold42 (.I(net56),
    .Z(net334));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold43 (.I(_01991_),
    .Z(net335));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold44 (.I(_00075_),
    .Z(net336));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold45 (.I(net386),
    .Z(net337));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold46 (.I(net86),
    .Z(net338));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold47 (.I(_02049_),
    .Z(net339));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold48 (.I(_00092_),
    .Z(net340));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold49 (.I(net389),
    .Z(net341));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold50 (.I(net58),
    .Z(net342));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold51 (.I(_02060_),
    .Z(net343));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold52 (.I(_00095_),
    .Z(net344));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold53 (.I(wbs_adr_i[22]),
    .Z(net345));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold54 (.I(net54),
    .Z(net346));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold55 (.I(net409),
    .Z(net347));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold56 (.I(_01995_),
    .Z(net348));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold57 (.I(_00076_),
    .Z(net349));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold58 (.I(net413),
    .Z(net350));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold59 (.I(net65),
    .Z(net351));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold60 (.I(net388),
    .Z(net352));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold61 (.I(net385),
    .Z(net353));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold62 (.I(net396),
    .Z(net354));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold63 (.I(net390),
    .Z(net355));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold64 (.I(wbs_adr_i[20]),
    .Z(net356));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold65 (.I(_01694_),
    .Z(net357));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold66 (.I(net384),
    .Z(net358));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold67 (.I(wbs_dat_i[12]),
    .Z(net359));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold68 (.I(net393),
    .Z(net360));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold69 (.I(net394),
    .Z(net361));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold70 (.I(net381),
    .Z(net362));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold71 (.I(net401),
    .Z(net363));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold72 (.I(net399),
    .Z(net364));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold73 (.I(net403),
    .Z(net365));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold74 (.I(net402),
    .Z(net366));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold75 (.I(net407),
    .Z(net367));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold76 (.I(net387),
    .Z(net368));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold77 (.I(net405),
    .Z(net369));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold78 (.I(net412),
    .Z(net370));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold79 (.I(net414),
    .Z(net371));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold80 (.I(_01746_),
    .Z(net372));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold81 (.I(net411),
    .Z(net373));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold82 (.I(net391),
    .Z(net374));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold83 (.I(net404),
    .Z(net375));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold84 (.I(net408),
    .Z(net376));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold85 (.I(wbs_cyc_i),
    .Z(net377));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold86 (.I(_01690_),
    .Z(net378));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold87 (.I(wbs_dat_i[6]),
    .Z(net381));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold88 (.I(wbs_dat_i[4]),
    .Z(net382));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold89 (.I(wbs_dat_i[10]),
    .Z(net383));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold90 (.I(wbs_dat_i[15]),
    .Z(net384));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold91 (.I(wbs_dat_i[19]),
    .Z(net385));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold92 (.I(wbs_dat_i[8]),
    .Z(net386));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold93 (.I(wbs_dat_i[29]),
    .Z(net387));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold94 (.I(wbs_dat_i[13]),
    .Z(net388));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold95 (.I(wbs_dat_i[11]),
    .Z(net389));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold96 (.I(wbs_dat_i[14]),
    .Z(net390));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold97 (.I(wbs_adr_i[21]),
    .Z(net391));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold98 (.I(_01987_),
    .Z(net392));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold99 (.I(wbs_dat_i[16]),
    .Z(net393));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(bus_in_gpios[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input10 (.I(bus_in_serial_ports[1]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input11 (.I(bus_in_serial_ports[2]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input12 (.I(bus_in_serial_ports[3]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(bus_in_serial_ports[4]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(bus_in_serial_ports[5]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(bus_in_serial_ports[6]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(bus_in_serial_ports[7]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(bus_in_timers[0]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(bus_in_timers[1]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input19 (.I(bus_in_timers[2]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(bus_in_gpios[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input20 (.I(bus_in_timers[3]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(bus_in_timers[4]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(bus_in_timers[5]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(bus_in_timers[6]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(bus_in_timers[7]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input25 (.I(io_in[0]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input26 (.I(io_in[10]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input27 (.I(io_in[11]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input28 (.I(io_in[12]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input29 (.I(io_in[4]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input3 (.I(bus_in_gpios[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input30 (.I(io_in[5]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input31 (.I(io_in[6]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input32 (.I(io_in[7]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input33 (.I(io_in[8]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input34 (.I(io_in[9]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(irqs[0]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input36 (.I(irqs[1]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input37 (.I(irqs[2]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input38 (.I(irqs[3]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input39 (.I(irqs[4]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input4 (.I(bus_in_gpios[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input40 (.I(irqs[5]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input41 (.I(irqs[6]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input42 (.I(rom_bus_in[0]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input43 (.I(rom_bus_in[1]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input44 (.I(rom_bus_in[2]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input45 (.I(rom_bus_in[3]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input46 (.I(rom_bus_in[4]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input47 (.I(rom_bus_in[5]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input48 (.I(rom_bus_in[6]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input49 (.I(rom_bus_in[7]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(bus_in_gpios[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input50 (.I(wb_rst_i),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input51 (.I(net371),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input52 (.I(net356),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input53 (.I(net374),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input54 (.I(net345),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input55 (.I(net377),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input56 (.I(net333),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input57 (.I(net329),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input58 (.I(net341),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input59 (.I(net307),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(bus_in_gpios[5]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input60 (.I(net352),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input61 (.I(net355),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input62 (.I(net358),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input63 (.I(net360),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input64 (.I(net361),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input65 (.I(net350),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input66 (.I(net353),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input67 (.I(net347),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input68 (.I(net354),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input69 (.I(net363),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(bus_in_gpios[6]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input70 (.I(net364),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input71 (.I(net365),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input72 (.I(net366),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input73 (.I(net369),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input74 (.I(net367),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input75 (.I(net375),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input76 (.I(net373),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input77 (.I(net368),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input78 (.I(net311),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input79 (.I(net376),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(bus_in_gpios[7]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input80 (.I(net370),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input81 (.I(net303),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input82 (.I(net315),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input83 (.I(net321),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input84 (.I(net362),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input85 (.I(net318),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input86 (.I(net337),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input87 (.I(net325),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input88 (.I(wbs_stb_i),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input89 (.I(wbs_we_i),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input9 (.I(bus_in_serial_ports[0]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap252 (.I(_01415_),
    .Z(net252));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output100 (.I(net100),
    .Z(RAM_end_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output101 (.I(net101),
    .Z(RAM_end_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output102 (.I(net102),
    .Z(RAM_end_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output103 (.I(net103),
    .Z(RAM_end_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output104 (.I(net104),
    .Z(RAM_end_addr[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output105 (.I(net105),
    .Z(RAM_end_addr[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output106 (.I(net106),
    .Z(RAM_start_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output107 (.I(net107),
    .Z(RAM_start_addr[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output108 (.I(net108),
    .Z(RAM_start_addr[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output109 (.I(net109),
    .Z(RAM_start_addr[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output110 (.I(net110),
    .Z(RAM_start_addr[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output111 (.I(net111),
    .Z(RAM_start_addr[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output112 (.I(net112),
    .Z(RAM_start_addr[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output113 (.I(net113),
    .Z(RAM_start_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output114 (.I(net114),
    .Z(RAM_start_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output115 (.I(net115),
    .Z(RAM_start_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output116 (.I(net116),
    .Z(RAM_start_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output117 (.I(net117),
    .Z(RAM_start_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output118 (.I(net118),
    .Z(RAM_start_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output119 (.I(net119),
    .Z(RAM_start_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output120 (.I(net120),
    .Z(RAM_start_addr[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output121 (.I(net121),
    .Z(RAM_start_addr[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output122 (.I(net122),
    .Z(WEb_raw));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output123 (.I(net123),
    .Z(boot_rom_en));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output124 (.I(net124),
    .Z(bus_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output125 (.I(net125),
    .Z(bus_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output126 (.I(net126),
    .Z(bus_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output127 (.I(net127),
    .Z(bus_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output128 (.I(net128),
    .Z(bus_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output129 (.I(net129),
    .Z(bus_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output130 (.I(net130),
    .Z(bus_cyc));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output131 (.I(net131),
    .Z(bus_data_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output132 (.I(net132),
    .Z(bus_data_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output133 (.I(net133),
    .Z(bus_data_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output134 (.I(net134),
    .Z(bus_data_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output135 (.I(net135),
    .Z(bus_data_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output136 (.I(net136),
    .Z(bus_data_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output137 (.I(net137),
    .Z(bus_data_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output138 (.I(net138),
    .Z(bus_data_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output139 (.I(net139),
    .Z(bus_we_gpios));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output140 (.I(net140),
    .Z(bus_we_serial_ports));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output141 (.I(net141),
    .Z(bus_we_timers));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output142 (.I(net142),
    .Z(cs_port[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output143 (.I(net143),
    .Z(cs_port[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output144 (.I(net144),
    .Z(cs_port[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output145 (.I(net145),
    .Z(io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output146 (.I(net146),
    .Z(io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output147 (.I(net251),
    .Z(io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output148 (.I(net148),
    .Z(io_oeb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output149 (.I(net149),
    .Z(io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output150 (.I(net150),
    .Z(io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output151 (.I(net151),
    .Z(io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output152 (.I(net152),
    .Z(io_oeb[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output153 (.I(net153),
    .Z(io_oeb[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output154 (.I(net154),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output155 (.I(net155),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output156 (.I(net156),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output157 (.I(net157),
    .Z(io_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output158 (.I(net158),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output159 (.I(net159),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output160 (.I(net160),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output161 (.I(net161),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output162 (.I(net162),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output163 (.I(net163),
    .Z(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output164 (.I(net253),
    .Z(io_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output165 (.I(net165),
    .Z(io_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output166 (.I(net166),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output167 (.I(net167),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output168 (.I(net168),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output169 (.I(net169),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output170 (.I(net170),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output171 (.I(net171),
    .Z(la_data_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output172 (.I(net172),
    .Z(la_data_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output173 (.I(net173),
    .Z(la_data_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output174 (.I(net174),
    .Z(la_data_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output175 (.I(net175),
    .Z(la_data_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output176 (.I(net176),
    .Z(la_data_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output177 (.I(net177),
    .Z(la_data_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output178 (.I(net178),
    .Z(la_data_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output179 (.I(net179),
    .Z(la_data_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output180 (.I(net180),
    .Z(la_data_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output181 (.I(net181),
    .Z(la_data_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output182 (.I(net182),
    .Z(la_data_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output183 (.I(net183),
    .Z(la_data_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output184 (.I(net184),
    .Z(la_data_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output185 (.I(net185),
    .Z(la_data_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output186 (.I(net186),
    .Z(la_data_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output187 (.I(net187),
    .Z(la_data_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output188 (.I(net188),
    .Z(la_data_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output189 (.I(net189),
    .Z(la_data_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output190 (.I(net190),
    .Z(la_data_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output191 (.I(net191),
    .Z(la_data_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output192 (.I(net192),
    .Z(la_data_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output193 (.I(net193),
    .Z(la_data_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output194 (.I(net194),
    .Z(la_data_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output195 (.I(net195),
    .Z(la_data_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output196 (.I(net196),
    .Z(la_data_out[32]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output197 (.I(net197),
    .Z(la_data_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output198 (.I(net198),
    .Z(la_data_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output199 (.I(net199),
    .Z(la_data_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output200 (.I(net200),
    .Z(la_data_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output201 (.I(net201),
    .Z(la_data_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output202 (.I(net202),
    .Z(la_data_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output203 (.I(net203),
    .Z(la_data_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output204 (.I(net204),
    .Z(le_hi_act));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output205 (.I(net205),
    .Z(le_lo_act));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output206 (.I(net206),
    .Z(reset_out));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output207 (.I(net207),
    .Z(rom_bus_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output208 (.I(net208),
    .Z(rom_bus_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output209 (.I(net209),
    .Z(rom_bus_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output210 (.I(net210),
    .Z(rom_bus_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output211 (.I(net211),
    .Z(rom_bus_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output212 (.I(net212),
    .Z(rom_bus_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output213 (.I(net213),
    .Z(rom_bus_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output214 (.I(net214),
    .Z(rom_bus_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output215 (.I(net215),
    .Z(wbs_ack_o));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output216 (.I(net216),
    .Z(wbs_dat_o[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output217 (.I(net217),
    .Z(wbs_dat_o[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output218 (.I(net218),
    .Z(wbs_dat_o[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output219 (.I(net219),
    .Z(wbs_dat_o[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output220 (.I(net220),
    .Z(wbs_dat_o[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output221 (.I(net221),
    .Z(wbs_dat_o[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output222 (.I(net222),
    .Z(wbs_dat_o[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output223 (.I(net223),
    .Z(wbs_dat_o[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output224 (.I(net224),
    .Z(wbs_dat_o[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output225 (.I(net225),
    .Z(wbs_dat_o[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output226 (.I(net226),
    .Z(wbs_dat_o[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output227 (.I(net227),
    .Z(wbs_dat_o[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output228 (.I(net228),
    .Z(wbs_dat_o[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output229 (.I(net229),
    .Z(wbs_dat_o[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output230 (.I(net230),
    .Z(wbs_dat_o[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output231 (.I(net231),
    .Z(wbs_dat_o[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output232 (.I(net232),
    .Z(wbs_dat_o[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output233 (.I(net233),
    .Z(wbs_dat_o[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output234 (.I(net234),
    .Z(wbs_dat_o[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output235 (.I(net235),
    .Z(wbs_dat_o[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output236 (.I(net236),
    .Z(wbs_dat_o[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output237 (.I(net237),
    .Z(wbs_dat_o[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output238 (.I(net238),
    .Z(wbs_dat_o[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output239 (.I(net239),
    .Z(wbs_dat_o[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output240 (.I(net240),
    .Z(wbs_dat_o[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output241 (.I(net241),
    .Z(wbs_dat_o[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output242 (.I(net242),
    .Z(wbs_dat_o[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output243 (.I(net243),
    .Z(wbs_dat_o[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output244 (.I(net244),
    .Z(wbs_dat_o[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output245 (.I(net245),
    .Z(wbs_dat_o[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output246 (.I(net246),
    .Z(wbs_dat_o[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output247 (.I(net247),
    .Z(wbs_dat_o[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output90 (.I(net90),
    .Z(RAM_end_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output91 (.I(net91),
    .Z(RAM_end_addr[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output92 (.I(net92),
    .Z(RAM_end_addr[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output93 (.I(net93),
    .Z(RAM_end_addr[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output94 (.I(net94),
    .Z(RAM_end_addr[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output95 (.I(net95),
    .Z(RAM_end_addr[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output96 (.I(net96),
    .Z(RAM_end_addr[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output97 (.I(net97),
    .Z(RAM_end_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output98 (.I(net98),
    .Z(RAM_end_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output99 (.I(net99),
    .Z(RAM_end_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer1 (.I(_00762_),
    .Z(net293));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer10 (.I(\as2650.cycle[3] ),
    .Z(net302));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer11 (.I(_00676_),
    .Z(net379));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer12 (.I(net379),
    .Z(net380));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer2 (.I(_01213_),
    .Z(net294));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer3 (.I(_00741_),
    .Z(net295));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer4 (.I(_01665_),
    .Z(net296));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer5 (.I(_00671_),
    .Z(net297));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer6 (.I(_00671_),
    .Z(net298));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 rebuffer7 (.I(_00794_),
    .Z(net299));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer8 (.I(_00752_),
    .Z(net300));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 rebuffer9 (.I(_00970_),
    .Z(net301));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire248 (.I(_02622_),
    .Z(net248));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_254 (.ZN(net254));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_255 (.ZN(net255));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_256 (.ZN(net256));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_257 (.ZN(net257));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_258 (.ZN(net258));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_259 (.ZN(net259));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_260 (.ZN(net260));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_261 (.ZN(net261));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_262 (.ZN(net262));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_263 (.ZN(net263));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_264 (.ZN(net264));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_265 (.ZN(net265));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_266 (.ZN(net266));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_267 (.ZN(net267));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_268 (.ZN(net268));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_269 (.ZN(net269));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_270 (.ZN(net270));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_271 (.ZN(net271));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_272 (.ZN(net272));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_273 (.ZN(net273));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_274 (.ZN(net274));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_275 (.Z(net275));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_276 (.Z(net276));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_277 (.Z(net277));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_278 (.Z(net278));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_279 (.Z(net279));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_280 (.Z(net280));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_281 (.Z(net281));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_282 (.Z(net282));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_283 (.Z(net283));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_284 (.Z(net284));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_285 (.Z(net285));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_286 (.Z(net286));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_287 (.Z(net287));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_288 (.Z(net288));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_289 (.Z(net289));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_290 (.Z(net290));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_291 (.Z(net291));
 assign io_oeb[0] = net275;
 assign io_oeb[13] = net256;
 assign io_oeb[14] = net257;
 assign io_oeb[15] = net258;
 assign io_oeb[16] = net259;
 assign io_oeb[17] = net260;
 assign io_oeb[18] = net261;
 assign io_oeb[1] = net254;
 assign io_oeb[2] = net255;
 assign io_oeb[4] = net276;
 assign io_out[0] = net262;
 assign io_out[4] = net263;
 assign irq[0] = net264;
 assign irq[1] = net265;
 assign irq[2] = net266;
 assign la_data_out[33] = net277;
 assign la_data_out[34] = net278;
 assign la_data_out[35] = net279;
 assign la_data_out[36] = net280;
 assign la_data_out[37] = net281;
 assign la_data_out[38] = net282;
 assign la_data_out[39] = net283;
 assign la_data_out[40] = net284;
 assign la_data_out[41] = net267;
 assign la_data_out[42] = net268;
 assign la_data_out[43] = net269;
 assign la_data_out[44] = net270;
 assign la_data_out[45] = net271;
 assign la_data_out[46] = net272;
 assign la_data_out[47] = net273;
 assign la_data_out[48] = net274;
 assign la_data_out[49] = net285;
 assign la_data_out[50] = net286;
 assign la_data_out[51] = net287;
 assign la_data_out[52] = net288;
 assign la_data_out[53] = net289;
 assign la_data_out[54] = net290;
 assign la_data_out[55] = net291;
endmodule

